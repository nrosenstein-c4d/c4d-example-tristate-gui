MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$       R�З������������������4����Ku���Ĉ-y�����Ks�����Kp�����Kq���čfq���čft���čfr����Rich���                PE  L ��R        � !  v  T      �^     �                                   @                   �� K   �� <                            � �                                   � @            � �                           .text   %t     v                   `.rdata  1   �  2   z             @  @.data   �   �     �             @  �.reloc  n   �     �             @  B                                                                                                                                                                                                                                                                                                                                                                                ��  �����������K  ������������L$t�   ù��  ������������  �����������j�h@fd�    P��V�P�3�P�D$ d�    �t$0���D$(    �9W  � �P�Qhdiem�B4�L$<�С �havem�@�L$8�@X�Ћ�L$Q���P@� ����QP���   havem�L$<�D$0�С ��L$���   Q� �D$, �Ѓ��D$4P���V  �L$4���D$(������%  �ƋL$ d�    Y^��$���������������j�hkfd�    P��(V�P�3�P�D$0d�    hTCAb�L$�^%  �L$�D$8    �-%  � ��t$D�@hdiem�@4�L$�D$@�ЋL$@�T$�R�T$R�P �L$���D$8 �K%  �L$�D$8�����:%  �ƋL$0d�    Y^��4�������̃�����V�B� �P����BPj?h�  �p~  j�D$P�F P���D$�  �D$    �~  �   ^������̸   �����������j�h�fd�    PQV�P�3�P�D$d�    �t$�L$�(  �L$�D$    ��t	�|.  ���3��L$�D$�����)  �ƋL$d�    Y^�����j�hgd�    P��$V�P�3�P�D$,d�    h�   j h���I h���A�  h�   h�  h��h� 舳  �� ��u�L$,d�    Y^��0á ��L$�@Q�@�С �j �@j��@�L$hؐQ�Ѓ��D$P�L$�D$8    �'  �L$�D$4��t�-  �L$���D$4 �(  ��L$�D$4 �(  3�� ��5l��@�L$�@Q�D$8�����С ��L$�@Q�@�С �j �@j��@�L$h�Q�Ѓ��D$P�L$�D$8   �&  �L$�D$4��t��,  �L$���D$4�(  ��L$�D$4�(  3�� ��5p��@�L$�@Q�D$8�����С ��L$�@Q�@�С �j �@j��@�L$h��Q�Ѓ��D$P�L$�D$8   ��%  �L$�D$4��t�T,  �L$���D$4�'  ��L$�D$4�t'  3�� ��5t��@�L$�@Q�D$8�����С ��L$�@Q�@�С �j �@j��@�L$h�Q�Ѓ��D$P�L$�D$8   �L%  �L$�D$4��t�+  �L$���D$4��&  ��L$�D$4��&  3�� ��5x��@�L$�@Q�D$8������jh(�h5  j��  �����t$�D$4   ��t���I  ���3�� ��L$�@Q�@�D$8�����С �j �@j��@�L$(hP�Q��V�D$4jP�D$T	   �&  � ����I�D$<�IP�D$X�����у�$�ƋL$,d�    Y^��0���hl��F/  hp��</  ht��2/  hx��(/  �������j�hCgd�    P��V�P�3�P�D$d�    ��t$�V�    �B    �D$$    ������D$    �D$    � �j ���   �L$�@QR�D$0�С ��L$���   Q� �D$4 �Ѓ��ƋL$d�    Y^�� ������������̡ ����   �AP���Y�����������̡ �Q���   � ��Y��������������̡ �Q�@�@��Y�髍  ������������t$�w  Y������V���x  �D$t	V�[  ����^� ��j�hhgd�    PQV�P�3�P�D$d�    ��t$�N �D$    �H;  ���D$�����)�  �D$t	V��  ���ƋL$d�    Y^��� ����V���;  �D$t	V��  ����^� ��j�h�gd�    PQVW�P�3�P�D$d�    ��jh0�h  j4��  �����|$�D$    ��tD���$  P�t$$���@�  �O �D$����]:  �G ���G�L$d�    Y_^��� 3��L$d�    Y_^��� ��������́|$�  V��u�����t$ ��  V�������   ^� ��̃��A �$�� R�T$R�D$    �P�$���������������j �� ��<  �����̃��A �T$�� R�T$R�D$    �P�$��������������QS�\$V�t$W�t$ �|$SW��V�D$�E  �L$h�  � ?  �t$ S�\$WV����B  �C��wv�$�x �=l���=p���=t���=x���tM� �W�@�@�Ћ �W�I���I�у���h   VPj j �5��5 ��5��5�W�B  _^[Y� �	   p  ���̋L$��t�j�� ���������������j�h�gd�    P��V�P�3�P�D$d�    �D$    �A0��u �L$,�����D$,�L$d�    Y^�� � �D$   �D$�t$,�D$$   �N�    �A    �    � �j ���   �T$�@RQ�D$0�Ћ ��D$���   P�	�D$   �D$4 �у��ƋL$d�    Y^�� � ������̸� ����������̡�� ��A�D$������A�D$��   � �D$� ��   � �������������̸D������������j�h(hd�    P��SUVW�P�3�P�D$,d�    ��� ��l$<�@j ���   hvdpi���Ћ �j �Qhacpi���   �͋��ҋ؁�suomt3��  � �3��@V���   hxvpi���ЉD$<� �V�@hyvpi���   ���ЉD$�D$P�D$@P���2C  K��   K�4  �L$��  h'  �\$8�  � ����QP�B8h�  �L$ ��h'  ��  � ����QP�B8h�  �L$ ��h'  ��  � ����QP�B8h�  �L$ �ЋGSjH�L$ Qh���h����p蛍  ��=�  |�����   ��S�ωW��8  �L$�   �D$4�����s  �Q�L$<��;�|S� �@�;�G�L$��;�|9��@�;�-�G@��   ��j �ωW�u8  �   h�  �w�C������ƋL$,d�    Y_^][��$� �������̋D$V�8��u�   �6W�x� �W���   �@8�Ѓ���w� �W���   �@8�Ѓ��3�_j �N �F0��7  �   ^� ̋ ��D$��t<�|$ �t$�I�t$�   t;�B�P���   �Ѓ�Ã�B�P���  �Ѓ�ù   ;�VB�W�xW�p�������u_^À|$ tWj V�= �������_�F��   ^�����������̋L$��t,�=� t�y���A�u
�D$�%t�� ��L$�@� �������������̋L$��t� ��L$�@��@  �����̡ �hﾭދ@��@  ��Y����������V�t$���t� �Q�@� �Ѓ��    ^�������������̡ ��@���  ���D$��t�x��u�   �3����������̡ ��@��  �� ��@��   ���D$�   ;�VB�W�xW�p�������u_^Ã|$ tWj V��; �������_�F��   ^���    �A    �A    �A    �����V��~ u=���t� �Q�@<�@�Ѓ��    W�~��t���{�  W�U������F    _^���������j�hXhd�    P��V�P�3�P�D$$d�    ��D$P� �  ��P���D$0    �-   �L$���D$,�����
�  �ƋL$$d�    Y^��(��������j�h�hd�    PQV�P�3�P�D$d�    ��~ uTjhP�j;j��������D$�D$    ��t�t$����  �3��D$�����F��u�L$d�    Y^��� �~ t3�9�"� ��t$�@<� �Ћȃ�3���F   �����L$d�    Y^��� ��������������V���F   � ��@<�@��3Ʌ����^��������������̋	� ���u�@� � �@<�t$�@Q�Ѓ�� ���������̃y t�   ËQ��u3�á �R�@<�1�@�Ѓ��������V��~ u=���t� �Q�@<�@�Ѓ��    W�~��t���[�  W�5������F    _^��������̋�� ���u�@� Ë@<�t$�@Q�Ѓ������������j�h�hd�    P��(SV�P�3�P�D$4d�    �D$    ����u� ��A�0�� ��t$H�@<Q�@�Ћ ������I�D$�IP�ѡ ��L$�@Q�@V�С ��L$0�@Q�@�D$L   �С �j �@j��@�L$<h��Q�Ѓ� � �j �@�L$�@@Q�L$,Q�L$ �D$H�Ѕ�� ��L$$�@Q�@���D$@�С ����@��tA�t$D�@V�Ћ ��D$�IP�I�D$   �D$D �у��ƋL$4d�    Y^[��4Ë@Hj�t$�L$�С �j��@j��t$T�@L�t$�L$$�С ��t$D�@V�@�С ��L$�@V�@Q�Ћ ��D$ �IP�I�D$    �D$L �у��ƋL$4d�    Y^[��4��j�hid�    P��(SV�P�3�P�D$4d�    �D$    ����u� ��A�0�� ��t$H�@<Q�@�Ћ ������I�D$�IP�ѡ ��L$�@Q�@V�С ��L$0�@Q�@�D$L   �С �j �@j��@�L$<h��Q�Ѓ� � �j �@�L$�@@Q�L$,Q�L$ �D$H�Ѕ�� ��L$$�@Q�@���D$@�С ����@��tA�t$D�@V�Ћ ��D$�IP�I�D$   �D$D �у��ƋL$4d�    Y^[��4Ë@Hj�t$�L$�С �j��@j��t$T�@L�t$�L$$�С ��L$$�@Q�@�С �j �@j��@�L$0h��Q�Ѓ�� �j �@�L$�@@Q�L$,Q�L$ �D$H�Ѕ�� ��L$$�@Q�@���D$@�С ����@��t�t$D�@V�������@Hj�t$�L$�С �j��@j��t$X�@L�t$�L$$�С ��t$D�@V�@�С ��L$�@V�@Q�Ћ ��D$ �IP�I�D$    �D$L �у��ƋL$4d�    Y^[��4����������j�hpid�    P��(SV�P�3�P�D$4d�    �D$    ����u� ��A�0�� ��t$H�@<Q�@�Ћ ������I�D$�IP�ѡ ��L$�@Q�@V�С ��L$0�@Q�@�D$L   �С �j �@j��@�L$<h��Q�Ѓ� � �j �@�L$�@@Q�L$,Q�L$ �D$H�Ѕ�� ��L$$�@Q�@���D$@�С ����@��tA�t$D�@V�Ћ ��D$�IP�I�D$   �D$D �у��ƋL$4d�    Y^[��4Ë@Hj�t$�L$�С �j��@j��t$T�@L�t$�L$$�С ��L$$�@Q�@�С �j �@j��@�L$0h��Q�Ѓ�� �j �@�L$�@@Q�L$,Q�L$ �D$H�Ѕ�� ��L$$�@Q�@���D$@�С ����@��t�t$D�@V�������@Hj�t$�L$�С �j��@j��t$X�@L�t$�L$$�С ��L$$�@Q�@�С �j �@j��@�L$0h��Q�Ѓ�� �j �@�L$�@@Q�L$,Q�L$ �D$H�Ѕ�� ��L$$�@Q�@���D$@�С ����@���D����@Hj�t$�L$�С �j��@j��t$\�@L�t$�L$$�С ��t$D�@V�@�С ��L$�@V�@Q�Ћ ��D$ �IP�I�D$    �\$L�у��ƋL$4d�    Y^[��4��������������j�h�id�    P��(SV�P�3�P�D$4d�    �D$    ����u� ��A�0�� ��t$H�@<Q�@�Ћ ������I�D$�IP�ѡ ��L$�@Q�@V�С ��L$0�@Q�@�D$L   �С �j �@j��@�L$<h��Q�Ѓ� � �j �@�L$�@@Q�L$,Q�L$ �D$H�Ѕ�� ��L$$�@Q�@���D$@�С ����@��tA�t$D�@V�Ћ ��D$�IP�I�D$   �D$D �у��ƋL$4d�    Y^[��4Ë@Hj�t$�L$�С �j��@j��t$T�@L�t$�L$$�С ��L$$�@Q�@�С �j �@j��@�L$0h��Q�Ѓ�� �j �@�L$�@@Q�L$,Q�L$ �D$H�Ѕ�� ��L$$�@Q�@���D$@�С ����@��t�t$D�@V�������@Hj�t$�L$�С �j��@j��t$X�@L�t$�L$$�С ��L$$�@Q�@�С �j �@j��@�L$0h��Q�Ѓ�� �j �@�L$�@@Q�L$,Q�L$ �D$H�Ѕ�� ��L$$�@Q�@���D$@�С ����@���D����@Hj�t$�L$�С �j��@j��t$\�@L�t$�L$$�С ��L$$�@Q�@�С �j �@j��@�L$0hĒQ�Ѓ�� �j �@�L$�@@Q�L$,Q�L$ �D$H�Ѕ�� ��L$$�@Q�@���D$@�С ����@��������@Hj�t$�L$�С �j��@j��t$`�@L�t$�L$$�С ��t$D�@V�@�С ��L$�@V�@Q�Ћ ��D$ �IP�I�D$    �\$L�у��ƋL$4d�    Y^[��4ËD$����EȉL$�(�  �������̡ ��@<�@����̋D$����u���VP�L$��  �D$P�D$P�L$�D$    �D$    �C�  ����   �t$��$    �D$��tB��t=��uZ� ��t$���   �@H�Ћ ��ЋA���@xV���Ѕ�u,�   ^��á ��t$���   �@T��VP�J�������uԍD$P�D$P�L$��  ���x���3�^����j�h!jd�    P��HSUVW�P�3�P�D$\d�    3ۉ\$� ��L$,�@Q�@�С �S�@j��@�L$8hȒQ�С ��L$@�@<Q�@�\$|�Ћ ����I�D$D�IPǄ$�   �����у���u3��L$\d�    Y_^][��T�V�L$(3���  �D$P�D$$P�L$,���  ���  �l$l���$    �|$ ��   � ��t$���   �@T�Ћ�����tc� ��D$<�IP�I�у��D$<Pj�D$T��P���D$p   �\$$�p  �Ћ ����AU�@x���D$h   �\$���D$��t�D$ �D$d   ��t� ��L$L�@����@Q�\$�Ѓ��D$d������t� ��L$<�@Q�@����Ѓ��|$ u�D$P�D$$P�L$,�ȿ  ��� �����|$�ǋL$\d�    Y_^][��T�����j�hvjd�    P��DSUVW�P�3�P�D$Xd�    �t$l3ۉ\$��u|� ��L$(�@Q�@�С �V�@j��@�L$4hԒQ�С ��L$<�@<Q�@�t$x�Ћ ����I�D$@�IP�D$|�����у���u3��L$Xd�    Y_^][��P�V�L$$3�蓾  �D$P�D$ P�L$(�о  ����   �|$h�d$ �D$����   � ��t$���   �@T�Ћ�����tc� ��D$8�IP�I�у��D$8Pj�D$P��P���D$l   �\$$�n  �Ћ ����AW�@x���D$d   �\$���D$l��t�D$l �D$`   ��t� ��L$H�@����@Q�\$�Ѓ��D$`������t� ��L$8�@Q�@����Ѓ��|$l tR�l$�ŋL$Xd�    Y_^][��PÃ�u3�L$��t+� �Q���   �@H�Ћ ��ЋA���@xW���Ѕ�t��D$P�D$ P�L$(�t�  �����������������̡ ��@<�@����̃=� uK����t� �Q�@<�@�Ѓ���    V�5���t����  V���������    ^������������j�h�jd�    P��VW�P�3�P�D$ d�    �t$8�D$    � ��t$8�@�T$���   R�Ћ�� ��|$0�IW�I�D$,   �ѡ �W�@V�@�Ћ ��D$�IP�I�D$   �D$8 �у��ǋL$ d�    Y_^�� � ������������������������̅�t�j������̡ ��@��  �� ��@��(  ��j�h�jd�    P�� �P�3�P�D$$d�    �D$    � ��T$�@R��   �ЋL$4P�D$0   ���  �L$�D$   �D$, �h�  �D$4�L$$d�    Y��,� �̡ ��@��$  �� ��@��  �� ��@���  �� ��@��  �� ��@���  �� ��@��x  �� ��@��|  �� ��@��d  �� ��@��p  �� ��@��t  ���D$V����t	V�z�������^� ̡ �V�@j �@j����Ћ�^��������̡ �V�@j �t$�@���Ћ�^� ���̡ �V�@�t$�@j����Ћ�^� ���̡ ��@�@����̡ �V�@j ���   ��L$j V�Ћ�^� �������������̡ ��t$�@Q�@�Ѓ�� �������̡ ��t$�@Q�@�Ѓ����@� ��̡ �h#  �t$�@�t$�@l��� ��̡ �hF  �t$�@�t$�@l��� ��̡ ��t$�@�@t�Ћ �P���   �@X�Ѓ�� ������̡ ��t$�@�@t�Ћ ��t$�Ћ��   R�@`�Ѓ�� ̡ ��t$�@���   �Ћȅ�u� � �Q���   �@�Ѓ�� �����������̡ ��@���   ��   � ��������� ������������̸   � �������̸   � �������̸   � �������̸   � ��������� �������������3�� �����������3�� �����������3�� �����������3�� ����������̸   � �������̸   � �������̸   � ��������3�� �����������3�� ����������̋L$�D$�A4�D$�A �D$��D$�A0�D$�A@5 �A8h< �A<m< �A@�= �AD�= �AHw< �ALr< �AP�< �Al�� �AX�< �A\�� �A`�� �Ad�� �AT|< �Ah�< �Ap�� �At�< �A(�A,    �����������́�   h�   �D$j P��! j ��$�   �D$��$�   ��$�   ��$�   P������$�   h�   �D$T�D$(P��$�   ��$�   j��  ���   �j�hVkd�    P��   SV�P�3�P��$�   d�    ����
  ����H  ��$�   �L$ �T�  � ��L$�@Q�@Ǆ$�       �С �j �@j��@�L$h�Q�Ѓ��D$P�L$<Ƅ$�   ��  ��$�   PƄ$�   �ޱ  �L$<QP�D$|PƄ$�   ��  �L$,QP�D$lPƄ$�   �Ζ  ���j j�PƄ$�   �  ���L$T��Ƅ$�   萑  �L$pƄ$�   ��  ��$�   Ƅ$�   �k�  �L$8Ƅ$�   �Z�  � ��L$�@Q�@Ƅ$�    �Ѓ��L$Ǆ$�   �����)�  ��t	V�	  ���Ƌ�$�   d�    Y^[�Ĩ   � V�t$���  �����^� ���������Q�J	  YË�`��`��`��`��`��` ��`(��`,��`@�����������3��������������̋D$�     3�� ̋�PP�   ���́��   V��$�   ��u
3�^���   �h�   �D$j P� ��$�   ���D$h�   �D$P��$�   ��Ήt$0�D$@5 �D$Pm< �D$T�= �D$X�= �D$\r< �D$`w< �PPj���  ��^���   �������j�t$��������uË��������`��`�����������̡ ��@��   �� �V�@�t$��$  �6�Ѓ��    ^��������������̡ �V�@��(  V�t$�Ѓ���^� ��������������̡ �Q�@�t$��,  �Ѓ�� ����̡ �Q�@�t$��,  �Ѓ����@� �D$��t�P�3ҡ �R�@Q��8  �Ѓ�� ��������̡ ��t$�@Q��<  �Ѓ�� ������t$� ��t$�@�t$��@  Q�Ѓ�� ������������̡ ��t$�@�t$��D  Q�Ѓ�� ̡ ��t$�@Q��H  �Ѓ�� �����j�h�kd�    P��VW�P�3�P�D$ d�    �t$4�D$    � �Q�@�L$��L  Q�Ћ�� ��|$<�IW�I�D$8   �ѡ �W�@V�@�Ћ ��D$(�IP�I�D$(   �D$D �у��ǋL$ d�    Y_^�� � ���̡ �Q�@��T  �Ѓ������������̡ �Q�@��P  �Ѓ������������̡ ��t$�@Q��X  �Ѓ�� ����̡ ��t$�@Q��l  �Ѓ�� ����̡ ��@��0  �� ��@��4  �� ��@��p  �� ��@��t  �� ��@��\  �� �V�@�t$��`  �6�Ѓ��    ^����������������t$� ��t$�@�t$��d  �t$�t$Q�Ѓ�� ������t$� ��t$�@�t$��h  �t$�t$Q�Ѓ�� ����̡ �Q�@�@�Ѓ�����������������t$� ��t$�@�t$�@X�t$Q�Ѓ�� �����������̡ ��t$�@Q�@\�Ѓ�� �������̡ �Q�@�@ ��Y�j�h�kd�    P��V�P�3�P�D$d�    � �h�  �@Q���   �L$Q��P� ��D$0    ���   �@8�Ћ ������   �D$�	P�D$4�����у��ƋL$d�    Y^����̡ ��@��   ���t$� ��t$�@�t$�@Q�Ѓ�� �t$� ��t$�@�t$���   �t$Q�Ѓ�� ��������̡ ��@�@$������t$� ��t$�@�t$�@(�t$Q�Ѓ�� �������������t$� ��t$�@�t$�@,�t$Q�Ѓ�� �������������t$$� ��t$$�@�t$$�@`�t$$�t$$�t$$�t$$�t$$�t$$Q�Ѓ�(�$ �������̡ �V�@W�@��W�Ћ �W�J���I���t$� ��t$�Q�t$�N�QHP�B4j j W�Ѓ�(_^� �t$� ��t$�@�t$�@4�t$�t$�t$�t$Q�Ѓ� � � ��t$�@�t$�@@Q�Ѓ�� ���̡ ��t$�@Q�@D�Ѓ�� �������̡ �Q�@�@L�Ѓ���������������̡ �Q�@�@L�Ѓ���������������̡ �Q�@�@P�Ѓ���������������̡ ��t$�@Q�@T�Ѓ�� �������̡ ��t$�@Q�@T�Ѓ�� �������̡ �Q�@�@h�Ѓ���������������̡ ��t$�@�t$���   Q�Ѓ�� �j�h ld�    P��V�P�3�P�D$d�    �t$4�D$    � ��t$4�@Q���   �L$Q�ЋЋt$<j �    �F    � �R���   V�@�D$@   �Ћ ��D$(���   P�	�D$(   �D$D �у� �ƋL$d�    Y^�� � �����������̡ ��@� �����̡ �V�@�t$�@�6�Ѓ��    ^���t$� ��t$�@�t$���   �t$�t$Q�Ѓ�� ����̡ �V�@�t$�@�6�Ѓ��    ^��QS�\$V�C    � ���@V�@h�Ѓ���� �u �@h����0  h�  �Ѓ�^3�[Y� �L$Q�L$Q�t$�D$    �@V���   �Ѓ���t�3�9t$~+W�d$ �D$�<� �<�tj����  ��t��F;t$|�_�D$P��������   ^[Y� ��QS�\$V�C    � ���@V�@h�Ѓ���� �u �@h����0  h�  �Ѓ�^3�[Y� �L$Q�L$Q�t$�D$    �@V���   �Ѓ���tσ|$ t�3�9t$~?W�D$����t+� �Q�@�@h�Ѓ���t�D$j�<�����
  ��t�8F;t$|�_�D$P��������   ^[Y� ������̡ ��@��x  �� ��@��|  �� �Q�@���   �Ѓ������������̡ ��t$�@Q���   �Ѓ�� ����̡ ��@���   �� �V�@�t$���   �6�Ѓ��    ^���������������VW���O��  W�f�G f�G(f�G0f�G8f�G@f�GHf�GPf�GX�    �G`    �Gd    �Gh    �Gp�Gx�����G|   ��_^�������j�h&ld�    PQV�P�3�P�D$d�    ��t$�D$    �k   �N�D$�����+�  �L$d�    Y^�������������W��    �A`    �Ad    �Ah    �Ap�Ax�����A|   ���������������SW�����t7��������xP t$V�������j j �pPj�GP�������H ���^�    �O`��t� �Q�@�@�Ѓ��G`    _[��������������j�h]ld�    PQ�P�3�P�D$d�    jh@�h�   h�   �i������D$�D$    ��t���/����L$d�    Y���3��L$d�    Y����������������j�h�ld�    PVW�P�3�P�D$d�    �|$�7��t,�t$���D$    ������N�D$����葂  V�k������    �L$d�    Y_^��á �S�@U�l$��   VW��W�_dS�wx�w`UV�Ѓ��G|����   �? ��   �; ��   �wpV�_hSU�
�  ����u&�W��� �h���@h  ��0  �Ѓ��wU���҆  �j j jV��  �G|��t��������G|_^][� �G|�Gx����_^][� �G|�����    � ��6�@�@�Ѓ��    �G|_^][� �����������V������W��    �F`    �Fd    �Fh    �Fp�Fx�����F|   ^������W���d �G`t~S�\$;_xtsU�/�͉D$�����xP u����%V���	���S�t$�pPj�GP��������H ���^�G|]��u�D$�_x��t�    �G`[_� �L$�Gx������t�3�[_� �̋D$��t	�Ap� �yd t�Ah� 3��y|��� ��������t$� ��t$�@�t$�@�t$�t$�t$�t$Q�Ѓ� � � ��t$�@Q�@�Ѓ�� �������̡ �Q�@�@��Yá ��t$�@�t$�@Q�Ѓ�� ���̡ ��@� �����̡ �V�@�t$�@�6�Ѓ��    ^��VW��������t$���t$�x@�t$�����H ���_^� �����VW�������t$���t$�xD�t$�����H ���_^� �����W���h����xH u3�_�V���V����ύpH�L����H �^_�����W���8����xL u3�_� V���$����t$���t$�pL�t$�����H ���^_� ��W��������xP u���_� V��������t$���t$�pP�t$�t$������H ���^_� �������������W�������xT u���_� V�������t$���t$�pT�����H ���^_� �����W���h����xX u���_� V���S����t$�ύpX�E����H ���^_� ���������j�h�ld�    P��$SVW�P�3�P�D$4d�    �ً|$D��tA�L$ �W������D$<    ������pL�D$ P��������H ��ЍL$ ��D$<���������t$H��tj� ��L$�@Q�@�С ��L$�@V�@Q�D$H   �С ��L$�@Q�@�D$L�����Ѓ����f����H@��t� �V�@Q�@�Ѓ��L$4d�    Y_^[��0� ��������VW���'����t$�΍xH�����H ���_^� �������������W��������x` u	� }  _� V��������t$�ύp`������H ���^_� �������SVW�������x` u� }  �$�������p`�D$���P�������H ��Ћ�� ��\$�IS�I�у�;�@� �S�@�@�Ѓ�;�+���O����t$���t$�pDS�t$�8����H ���_^[� _^�����[� W�������xP u	�����_� V�������t$ ���t$ �pP�t$ �t$ �t$ �t$ ������H ���^_� ���W��������xT u	�����_� V�������t$���t$�pT�����H ���^_� ���W�������xX tV���z����t$�ύpX�l����H ���^_� ���$P�t$ �D$    �D$    �D$    �D$    �D$    �D$    ���  ����t,�$��t%�t$� ��t$�@�t$�@X�t$Q�Ѓ����3�������������z  �����������SUV��L$�F�.�V���    �;�~|�
W�@�+����ρ�  �yI���Au��u	�   +��� �h0��Hh�   ��    P��  U�ЋЃ���t�N�~_�^�^]��[� �F_�F^]��[� �^^][� ��������������A    �A    �A    �����V��~ ���u� ��v�@4� �Ѓ��F    �F    ^���������������̸   ����������̸   �����������3�� ������������ ������������̡ �V�@4��@$h�  �v���t$� ��t$�@4�t$�@�t$�v�Ѓ�2�^� ����������������t$��t$�t$�t$�P� ��������3�� ����������̸   � ��������� �������������Q� �U�@V�@ W�|$���3���=INIb�!  �  =SACbqt(=$'  t
=MicM�i  �E W���P$�   _��^]Y� �E �L$Q�L$Q�͉t$�t$�P��t�t$� ��t$�@4�u�@�Ѓ��   _��^]Y� =ARDb�  � �S�@j ���   j���Ћء �j �@j���   ���ЋL$��� �j �@j���   �ЋL$�� �j �@j���   ���t$�U PVWS���R[�   _��^]Y� �E ���P�   _��^]Y� =NIVb\tD=NPIbt-=ISIbuS�u ����  P���  P���V�   _��^]Y� �E W���P_^]Y� �E ���P�   _��^]Y� =cnyst	_��^]Y� � �j �@hIicM���   ���ЋU WP���R _^]Y� ������������j�h�ld�    P��,V�P�3�P�D$4d�    ��~ ��   � ��v�@4�@�Ѓ|$H t+� �P�F�I0�p�Al�Ѓ��L$4d�    Y^��8� ���L$ hARDb�D$�D$    ������NP�D$P�D$P�D$H    �  � ��L$���   Q� �Ѓ��L$ �D$<����������L$4d�    Y^��8� ����������̡ ��t$�@4�q�@l�Ѓ��   � ̡ ��q�@4�@�Ѓ�������������̡ ��q�@4�@�Ѓ�������������̡ ��q�@4�@�Ѓ�������������̡ ��q�@4�@|�Ѓ�������������̡ ��q�@4���   �Ѓ����������̡ ��t$�@4�q�@(�Ѓ�� �������t$� ��t$�@4�t$�@,�q�Ѓ�� ���������������t$� ��t$�@4�q�@0�Ѓ�� �̡ ��q�@4�@4��Y��������������̡ ��t$�@4�q���   �Ѓ�� ��̡ ��t$�@4�q�@ �Ѓ�� �����̡ ��t$�@4�q�@$�Ѓ�� �����̡ �V���   �t$�@WV���Ѓ���� �V���   u�@@�Ћ �P�I4�w�A �Ѓ�_^� �@�Ѓ���� �u&���   V�@8�Ћ �P�I4�w�A$�Ѓ�_^� �@h���0  h
  �Ѓ�_^� ����������������t$� ��t$�@4�q�@D�Ѓ�� ���t$� ��t$�@4�q�@H�Ѓ�� ���t$� ��t$�@4�q�@L�Ѓ�� ���t$� ��t$�@4�q�@P�Ѓ�� �̡ �S���   V�@W�|$W���Ѓ���� ����   �@��   �t$V�Ѓ���� �V���   u5�@@�Ћ �W���   ���I@�ы �V�I4P�s�AP�Ѓ�_^[� �@�Ѓ���� �u<���   V�@8�Ћ �W���   ���I@�ы �V�I4P�s�AH�Ѓ�_^[� �@h,���0  h�  �Ѓ�_^[� W�Ѓ���� ���   ���   �t$�@V�Ѓ���� �V���   u5�@@�Ћ �W���   ���I8�ы �V�I4P�s�AL�Ѓ�_^[� �@�Ѓ���� �u<���   V�@8�Ћ �W���   ���I8�ы �V�I4P�s�AD�Ѓ�_^[� �@hL���0  h�  �Ѓ�_^[� �@hl���0  h�  �Ѓ�_^[� ����������t$� ��t$�@0�t$���   �t$�q�Ѓ�� ������̡ ��t$�@0�q���   �Ѓ�� ����D$� ����@0�$�t$���   �t$�q�Ѓ�� ��t$� ��t$�@4�t$�@�t$�q�Ѓ�� �����������t$� ��t$�@4�t$�@�t$�q�Ѓ�� �����������t$(� ��t$(�@4�t$(�@T�t$(�t$(�t$(�t$(�t$(�t$(�t$(�q�Ѓ�,�( ���t$� ��t$�@4�t$��  �t$�q�Ѓ�� ��������t$ �D$�t$ � ��t$ �@4�t$ ��  ���D$�D$$�$�q�Ѓ�$�  ������������̡ �h�����@4h�����@Th�����t$�t$h����h����h����h�����t$(�q�Ѓ�,� ����������̡ ��t$�@4�q�@8�Ѓ�� �����̡ ��t$�@4�q�@<�Ѓ�� �������t$� ��t$�@4�q���   �Ѓ�� ��������������̡ ��q�@4�@@�Ѓ�������������̡ ��q�@4��  �Ѓ����������̡ ��D$�@4����  �$�q�Ѓ�� ����������t$� ��t$�@4�t$�@X�t$�q�Ѓ�� ���������̡ ��q�@4�@`��Y��������������̡ ��q�@4�@d�Ѓ���������������t$� ��t$�@4�t$��   �t$�q�Ѓ�� ��������t$� ��t$�@4�t$�@\�t$�t$�t$�q�Ѓ�� ���t$� ��t$�@4�q��  �Ѓ�� ����������������t$� ��t$�@4�q�@h�Ѓ�� ���t$� ��t$�@4�q��  �Ѓ�� ����������������t$� ��t$�@4�q�@p�Ѓ�� ��j�h�ld�    P��VW�P�3�P�D$ d�    ��hYALf�L$�;���P� ��w�B4�D$0    �@l�Ѓ��L$�D$(�����M����L$ d�    Y_^�� ������������UVW�|$���t� ��L$�@j ���   j�Љ�t$��t� ��L$�@j ���   j�Љ� �V�@4W�u�@p�Ѓ�_^]� �������������t$� ��t$�I�@0�t$���   �q�Ѓ�� ���������t$� ��t$�@4�t$�@x�t$�q�Ѓ�� ���������̡ ��t$�@4�q�@t�Ѓ�� �������t$� ��t$�@4�t$���   �t$�t$�q�Ѓ�� ����t$� ��t$�@4�t$���   �t$�t$�q�Ѓ�� ��̃�� �SW�D$    �D$    �@�ًL$$���   �{j j�ЋL$$�D$� �j �@j���   �ЉD$� ��L$�@0Q�@`�L$Q�w�С ��s�@4�@�Ћ �j �I0�T$,R�T$4R�T$(R�T$4RP�C�p�Ah�Ѓ�,�|$( _[t.�|$$ t.�L$�T$;�~C�D$�;�}9�$�T$;�~.�D$��|$$ u�L$�T$;�~�D$�;�}�   ��� 3���� ����������������t$�D$� ����@4�D$�D$���   �$�t$�q�Ѓ�� ������t$� ��t$�@4�t$���   �q�Ѓ�� ����������̡ ��q�@4���   �Ѓ����������̡ ��q�@4��  �Ѓ�����������V��V��� �h�� �@0� �Ѓ��F�F    ��^�����V��N����t� �Q�@0�@�Ѓ��F    ^������̸   ����������̸   ����������̸   � ��������3�� �����������3���������������� ����������������������������̡ �V�@W�|$�@ �����=NIVb��   ��   =TCAbttK=$'  t2=MicM��   � �j �@hIicM���   ���ЋWP���R_^� �W���P_�   ^� � �j �@hdiem���   ���ЋWP���R_^� =INIbuz�~ u���F   �P_^� �~ t�����P_^� =atni=t/=ckhct=ytsdu8����P_�F    3�^� ����P_^� �N�  _3�^� =cnys����_3�^� �����V��N��u3�^� � �j �@0j ���   j j j �t$4j �t$(jQ���t$D� ��t$D�@0�t$D���   �t$Dj �t$D�v�Ѓ�D^� ��������̋I��u3�á �Q�@0�@�Ѓ�����̋I��u3�� � �Q�@0�@�Ѓ�� j�h7md�    P��V�P�3�P�D$d�    �D$    �q��u �D$,�    �p�L$d�    Y^�� � �D$0�H�� �Q�t$8�@0R���   �L$VQ�ЋЋt$@j �    �F    � �R���   V�@�D$D   �Ћ ��D$,���   P�	�D$,   �D$H �у�$�ƋL$d�    Y^�� � �������������̡ ��t$�@0�q���   �Ѓ�� ��̡ ��q�@0���   �Ѓ����������̡ �j �@0j ���   j j j j j j j4�q�Ѓ�(�������̡ �j �@0j ���   j j j j j j j;�q�Ѓ�(�������̡ ��t$�@0�q�@�Ѓ�� �����̋I��t(� �j �@0j ���   j j j j �t$j jQ�Ѓ�(� ���������������t$� ��t$�@4�t$�@,�q�Ѓ�� ���������������t$� ��t$�@4�q�@0�Ѓ�� �̡ ��q�@4�@4��Y���������������V�q��u3�^� �D$�H�� �Q�t$�@0R�@V�Ѓ�^� ��������������V�q��u3�^� �D$�H�� �Q�@0R���   V�Ѓ�^� ��������������̋D$3�h�����h  ���Pj BRj �t$ �t$ �   � ����j�hbmd�    P��$VW�P�3�P�D$0d�    ��htniv�L$ ������ ��t$D�@hulav�@4�L$$�D$@    �С �hgnlf�@htmrf�@4�L$$�С ��t$H�@hinim�@4�L$$�С ��t$L�@hixam�@4�L$$�С ��t$P�@hpets�@4�L$$�С ��t$T�@hsirt�@4�L$$�ЋL$X�t$\��  �u�����t.� �Q�@h2nim�@4�L$$�С �V�@h2xam�@4�L$$�ЍD$P�t$D�D$P������P� ��D$<���   �@8�Ћ ������   �D$�	P�D$@ �у��L$�D$8����������ƋL$0d�    Y_^��0�  ��������������U����j�h�md�    P��pV�P�3�P�D$xd�    ��htlfv�L$4�6���� ��E�@���@,�$hulav�L$<Ǆ$�       �С ��u,�@htmrf�@4�L$8�С ��E�@���@,�$hinim�L$<�С ��E�@���@,�$hixam�L$<�С ��E$�@���@,�$hpets�L$<�С ��uD�@hsirt�@4�L$8���U0W�f.џ��Dz�E8f.����D{A� ����@�$�@,h2nim�L$<�С ��E8�@���@,�$h2xam�L$<�С ��u@�@hdauq�@4�L$8�ЍD$0P�u�D$$P������P� �Ƅ$�   ���   �@8�Ћ ������   �D$ �	PƄ$�    �у��L$0Ǆ$�   ����������ƋL$xd�    Y^��]�@ ����������t$(W�j ���D$�$�D$8htemf�� �D$�D$T�D$�D$L�D$�D$D�$�t$@�����( �������L$f.������%Ж���D{�Y��^��T$f.����D{�Y��^��t$(W�j ���D$�$�D$8�Y�hrgdf�� �^��D$�D$D�L$�T$�$�t$@�����( ���t$(�ȖW�j ���D$�$�D$8�^�htcpf�� �D$�D$T�^��D$�D$L�^��D$�D$D�$�t$@�����( ��U����j�h�md�    P��hSVW�P�3�P�D$xd�    �ًE��u)� ��@���   �Ѕ�u�L$xd�    Y_^[��]� �����  htlfv�L$4�������ufn�������YǄ$�       �D$�D$�$��  �F�\$$�D$�D$�$�q�  �D$$�\$�^D$� ��$�@hulav�@,�L$<�С �hmrff�@htmrf�@4�L$8�Ћufn�������Y�D$$�D$$�$��  �F�\$�D$$�D$$�$���  �D$�\$$�^D$$� ��$�@hinim�@,�L$<�Ћufn�������Y�D$$�D$$�$��  �F�\$�D$$�D$$�$��  �\$$�D$�^D$$� ��$�@hixam�@,�L$<�С �����@���@,�$hpets�L$<�С �j �@hdauq�@4�L$8�С �W�@hspff�@4�L$8�С ��u �@hsirt�@4�L$8�ЍD$0P�u�D$$P������P� �Ƅ$�   ���   �@8�Ћ ������   �D$ �	PƄ$�    �у��L$0Ǆ$�   ���������ƋL$xd�    Y_^[��]� ��������������j�h�md�    P��$V�P�3�P�D$,d�    ��hCITb�L$������ ��t$@�@hCITb�@8�L$ �D$<    �С ��t$D�@hsirt�@4�L$ �С ��t$H�@hulav�@4�L$ �ЍD$P�t$@�D$P���q���P� ��D$8���   �@8�Ћ ������   �D$�	P�D$< �у��L$�D$4���������ƋL$,d�    Y^��0� �����V�q��u3�^� �D$�D$�H�� �Q�t$$�@0���@(�D$�D$(�$�t$$RV�Ѓ�$^� j�hnd�    P��V�P�3�P�D$d�    ��L$,�D$P��Z  j �t$4��P�t$4�D$0    �b���� ����I�D$�IP�D$$�����у��ƋL$d�    Y^��� �������������V�q��u3�^� �D$�H�� �Q�@0�L$�@,QRV�ЋL$3҃�9T$^�� ��������������V�q��u3�^� �D$�H�� �Q�t$�@0R�@,V�Ѓ�^� ��������������V�q��u3�^� �D$�H�� �Q�t$�@0R�@0V�Ѓ�^� ��������������UVW���O����   �D$�l$�P�0� �R�@0U�@0VQ�Ѓ���tb� t\�D$�H�� �Q�p0�EP�F0R�w�Ѓ���t6���t/�D$�H�� �Q�p0�EP�F0RW�Ѓ���t_^�   ]� _^3�]� �QV�q��u3�^Y� �D$W�H�� �Q�L$�D$    �@0Q�@8RV�Ћ�����t=�T$��t5� ��t$�AR�@�Ћt$����t� �V�@�@��V趩������_^Y� �����������V�q��u3�^� �D$�H�� �Q�t$�@0�t$�@<RV�Ѓ�^� ���������̋D$��V���u� ��@���   �Ѕ�u^��� W���?�  �v����t#�D$$�H�� �Q�@0�L$�@0QRV�Ѓ���fn�������Yؖ�L$ �D$�D$�Yؖ�$�.�  �~ �L$,_f��~@��f�A^��� ��������������j�h)nd�    P��V�P�3�P�D$d�    �� ��L$�@Q�@�Ѓ��D$P�t$,���D$(    ��������t�L$,�D$P��W  � ��D$�IP�I�D$$�����у��ƋL$d�    Y^��� ������V�q��u3�^� �D$�H�� �Q�@0j ���   j j j j j Rj1V�Ѓ�(^� ̡ �V�@j �t$���   ��L$��h���h  �j j jj P�t$$���%���^� ̡ �V�@j �t$���   ��L$���t$$���t$$j �t$(�t$(�t$(P�t$$�����^�  �������������U������<� �V�@�����   W��$�u��M���\$8�E8j �u@�΃��D$�E0�$�u,�E$�� �D$�E�D$�E�D$�D$t�$�u�����^��]�< ���������������U������<� �V�@�����   W��$�u��M���\$8j j ��W��D$�$�E$htemf�� ���D$�E�D$�E�D$�D$t�$�u�L���^��]�$ �����U������<� �V�@�����   W��$�u��M���\$8�Uf.������%Ж���D{�Y��^��Mf.����D{�Y��^�j j ��W��D$�$�E$�Y�hrgdf�� ���^��D$�D$t�T$�L$�$�u�x���^��]�$ �U������<� �V�@�����   W��$�u��M���\$8�Ȗj W�j �����D$�$�E$�^�htcpf�� �D$�E�^��D$�E�^��D$�D$t�$�u�����^��]�$ ̃�0� �V��W��D$����L$Q�t$H�D$�@�L$,���   Q�L$L���~ j �t$Tf�D$�t$T�~@�t$T�D$$P�t$P���t$Pf�D$8�����^��0� ���j�hTnd�    P�� V�P�3�P�D$(d�    �� ��L$�@Q�@�Ѓ��L$<�D$P�t$D�D$ P�D$<    �����t$D��j P�t$D�D$@����� ����I�D$�IP�D$4 �ѡ ��L$�@Q�@�D$8�����Ѓ��ƋL$(d�    Y^��,� ���j�h�nd�    P��HV�P�3�P�D$Pd�    ��L$4�QO  �L$dP�t$l�D$ P�D$d    �VI  �L$Q���D$\��Q  j j P�t$l���D$h�`���� ����I�D$�IP�D$\�у��L$�D$X ��P  �L$4�D$X������P  �ƋL$Pd�    Y^��T� ���������������U������x�U���V�uW���D$0���t.� ����@W����   �$R�����\$0�D$0�D$0� �W��L$8Q�u�D$@�D$H�D$P�@�L$p���   Q�����~ �wf�D$P�~@f�D$X�~@f�D$`��u
3�_^��]� �E�E�H�� �Q�u �@0���@(�D$�D$H�$�L$hQRV�Ѓ�$_^��]� ���V�q3���t,�D$�H�� �Q�@0�L$�@,QRV�Ћ�3���9D$��� �P�Q�t$�L$�R0�ҋ�^� �������������V�q��t#�D$�H�� �Q�@0�L$�@,QRV�Ѓ���� ��t$�A�t$�L$�@4�Ћ�^� ����̃�V�q��t#�D$�H�� �Q�@0�L$�@0QRV�Ѓ���� ��D$�A�L$�@,���$�t$ �Ћ�^��� ����̃�V�D$P�t$ W��t$ �D$����D$������ ����Q�L$ �R@�D$P�t$(�ҋ�^��� ������������̃�V��W�~W��D$�D$�D$����   �D$$�H�� �Q�@0�L$�@0QRW�Ѓ���t�~��tx�D$(�H�� �Q�@0�L$�@0QRW�Ѓ���tS�v��tL�D$,�H�� �Q�@0�L$�@0QRV�Ѓ���t'� ��L$�@Q�t$8�L$8�@H��_�   ^��� _3�^��� �����������j�h�nd�    P��V�P�3�P�D$d�    �� ��L$�@Q�@�Ѓ��D$P�t$,���D$(    ����� ����Q�L$,�R8�D$P�t$4�ҡ ��L$�@Q�@�D$$�����Ѓ��ƋL$d�    Y^��� ��������������j�h�nd�    P��V�P�3�P�D$$d�    ��L$�J  �D$P�t$8���D$4    ����� ����Q�L$8�R<�D$P�t$@�ҍL$�D$,�����+L  �ƋL$$d�    Y^��(� �����̃� V�qW��D$�D$�D$��t(�D$(�H�� �Q�@0�L$�@<Q�L$QRV�Ѓ����T$0���t� ��A�L$�@HQ�L$0R�ЋT$4���t � ��D$�@�L$,�@,���$R�Ћ�^�� � ����̋D$3҃8V�p�¸   h���h  ���E�3�����Rj @Pj V�t$$����^� �T$�t$3��:�t$��P�t$ �t$ �t$ �r�t$ ����� �T$�D$03��:��P�t$<���D$�D$@�$�t$<�D$8�� �D$�D$P�D$�D$H�D$�B�$�t$@�����8 ���̋D$3҃8�H��W�Rj ���D$�$�D$4htemf�� �D$�D$P�D$�D$H�D$�$�t$@�Q����  �������������̋D$�T$�h����%Ж3҃8��f.�����D{�Y��^��L$f.����D{�Y��^�Rj ��W��D$�$�D$4�Y�hrgdf�� �^��D$�T$�L$�,$�t$@�����  ���������̋D$�Ȗ3҃8W����PRj ���D$�$�D$4�^�htcpf�� �D$�D$P�^��D$�D$H�^��D$�$�t$@�����  ���������̋T$3��:��P�t$�B�t$�t$P�t$�t$�V���� ��̋D$�t$3҃8��RP�t$����� ���������������j�hod�    P��$V�P�3�P�D$,d�    ��hgnrs�L$�����D$@�D$4    �D$   �D$� ��L$�@Q���   j�L$ �D$<�С ��L$���   Q� �D$8 �ЋD$H���D$   �D$� ��L$�@Q���   j�L$ �D$<�С ��L$���   Q� �D$8 �Ѓ��D$P�t$@�D$P������P� ��D$8���   �@8�Ћ ������   �D$�	P�D$< �у��L$�D$4�����0����ƋL$,d�    Y^��0� �����������W�y��u3�_� �D$�D$�H�� �V�p0�D$Q�t$(�����D$�D$,�$P�F(RW�Ѓ�$^_� ���������̡ �j �@0j ���   j j j j j j j �q�Ѓ�(�������̋I��u3�� � ��t$�@4�t$��  Q�Ѓ�� ����̋I��u3�� � ��t$�@4�t$�@hQ�Ѓ�� �������̋I��u3�� � ��t$�@4�t$�@pQ�Ѓ�� �������̋I��u3�� � ��t$�@4�t$��  Q�Ѓ�� ������t$� ��t$�@0�t$���   �t$�q�Ѓ�� ������̡ ��P0�D$�pj j j �t$�t$j �0���   j=�q�Ѓ�(� �����������̡ ��P0�D$�p�t$j j j��t$j �0���   j=�q�Ѓ�(� �����������̋D$�t$����EС ��2�@0�t$�@@�q�Ѓ�� ��Q�I��u3�Y� � ��$Rj j �t$ �D$    �t$ �@0�t$ ���   �t$0�t$$jQ�ЋD$(��(Y� Q�I��u3�Y� � ��$Rj j �t$ �D$    �t$ �@0�t$ ���   �t$0�t$$jQ�ЋD$(��(Y� Q�I��u3�Y� � ��$Rj �t$$�D$    �t$ �@0�t$ ���   �t$ �t$0�t$$jQ�ЋD$(��(Y� ��������������Q�I��u3�Y� � ��$Rj �t$ �D$    �t$ �@0�t$ ���   �t$ j �t$$jQ�ЋD$(��(Y� Q�I��u3�Y� � ��$Rj �t$ �D$    �t$ �@0�t$ ���   �t$ j �t$$jQ�ЋD$(��(Y� Q�I��u3�Y� � ��$Rj �t$ �D$    �t$ �@0�t$ ���   �t$ j �t$$j*Q�ЋD$(��(Y� Q�I��u3�Y� � ��$Rj j �t$ �D$    �t$ �@0�t$ ���   j �t$$jQ�ЋD$(��(Y� ��Q�I��u3�Y� � ��$Rj j �t$ �D$    �t$ �@0�t$ ���   j �t$$jQ�ЋD$(��(Y� ��Q�I��u3�Y� � ��$Rj j �t$ �D$    �t$ �@0�t$ ���   j �t$$j	Q�ЋD$(��(Y� ��Q�I��u3�Y� � ��$Rj j �t$ �D$    �t$ �@0�t$ ���   j �t$$j
Q�ЋD$(��(Y� ��Q�I��u3�Y� � ��$Rj �t$ �D$    �t$ �@0�t$ ���   �t$ j �t$$jQ�ЋD$(��(Y� Q�I��u3�Y� � ��$Rj �t$ �D$    �t$ �@0�t$ ���   �t$ j �t$$jQ�ЋD$(��(Y� Q�I��u3�Y� � ��$Rj j �t$ �D$    �t$ �@0�t$ ���   �t$0�t$$j'Q�ЋD$(��(Y� Q�I��u3�Y� � ��$Rj j �t$ �D$    �t$ �@0�t$ ���   �t$0�t$$j,Q�ЋD$(��(Y� Q�I��u3�Y� � ��$Rj �t$ �D$    �t$ �@0�t$ ���   �t$ j �t$$j:Q�ЋD$(��(Y� Q�I��u3�Y� � ��$Rj j j �t$�D$    �t$ �@0j ���   j j)Q�ЋD$(��(Y� ������Q�I��u3�Y� � ��$Rj j �t$�D$    �@0j �t$ ���   j j j)Q�ЋD$(��(Y� �����̋I��u3�� � �j �@0j ���   j �t$�t$�t$j �t$ jQ�Ѓ�(� ���Q�I��u3�Y� � ��$Rj �t$ �D$    �t$ �@0�t$ ���   �t$ j �t$$jQ�ЋD$(��(Y� Q�I��u3�Y� � ��$Rj �t$ �D$    �t$ �@0�t$ ���   �t$ j �t$$j>Q�ЋD$(��(Y� Q�I��u3�Y� � ��$Rj j �t$ �D$    �t$ �@0�t$ ���   j �t$$jQ�ЋD$(��(Y� �̡ �j �@0j ���   j �t$�t$�t$j �t$ j.�q�Ѓ�(� �������������V�q��u3�^� �D$�H�� �Q�@0j ���   j j j �t$ �t$(RjV�Ѓ�(^� �������������V�q��u3�^� �D$�H�� �Q�@0j ���   j j j j j RjV�Ѓ�(^� �V�q��u3�^� �D$�H�� �Q�t$�@0R�@\V�Ѓ�^� �������������̃�SVW�t$ �ٍL$�+a  �D$ P�D$P�L$�ha  ��tm�|$�L$ ��tJ� �Q���   �@H�ЋS������tR�w� �j �A0j ���   j j �t$ V�7jR�Ѓ�(��t%�D$ P�D$P�L$��`  ��u�_^�   [��� _^3�[��� ��������������Q�I��u3�Y� � ��$Rj j �t$ �D$    �t$ �@0�t$ ���   j �t$$jQ�ЋD$(��(Y� �̡ �V�@4W�|$� �w���ЋD$�G    �w�H�� �Q�t$�@0W���   R�v�Ѓ�3Ʌ����G_^��� �������̋I��u3�� � �j �@0j ���   j �t$�t$�t$j �t$ j/Q�Ѓ�(� ��̋T$��u3�� �r�B    � ��t$�@0�q���   �Ѓ�� �����������̋I��u3�� � �j �@0j ���   j j j �t$j j jQ�Ѓ�(� ��������̡ �j �@0j ���   j j j j j j j6�q�Ѓ�(�������̋I��u3�� �t$� ��t$�@0�t$�@DQ�Ѓ�� ���̋I��u3��  �t$ � ��t$ �@0�t$ ���   �t$ �t$ �t$ �t$ �t$ Q�Ѓ�$�  ������������̋I��u3�á �Q�@0�@X�Ѓ�����̋I��u3�� � ��t$�@0�t$�@LQ�Ѓ�� �������̋Q��u3�� � ��H0�D$   �P�APR�Ѓ�� �����̋I��u3�� � ��t$�@0Q�@P�Ѓ�� �����������̋I��u3�� �t$� ��t$�@0�t$�@T�t$Q�Ѓ�� j�h+od�    P��VW�P�3�P�D$ d�    ���L$�����D$0�L$�P�0� �R�@0Q���   j j j j j Vj8�w�D$P    �Ћ���(��t�L$4�D$P�����L$�D$(���������ƋL$ d�    Y_^�� � ����������̋D$V�P�0� �R�t$�@0j ���   j j j j Vj9�q�Ѓ�(^� ���������̋D$V�P�0� �R�t$�@0�t$�@h�t$�t$V�q�Ѓ�^� �������������UVW�|$���t� ��L$�@j ���   j�Љ�t$��t� ��L$�@j ���   j�Љ� �V�@0W�u�@`�Ѓ�_^]� �������������t$� ��t$�@0�t$���   �q�Ѓ�� ����������̋T$� ��@0��t*���   R�q�Ћ ��t$�ЋA0R���   �Ѓ�� �t$�@|�q�Ѓ�� �����t$� ��t$�@0�t$�@p�t$�t$�q�Ѓ�� �������t$� ��t$�@0�t$�@d�t$�t$�q�Ѓ�� �����̡ �j �@0j �t$���   �t$ �t$ �t$j �t$ j3�q�Ѓ�(� ����������̋D$j �� �j �@0j ���   j j j j Rj�q�Ѓ�(� �D$j �� �j �@0j ���   j j jj Rj�q�Ѓ�(� �D$j �� �j �@0j ���   j j j j Rj�q�Ѓ�(� �D$V�P�0� �R�@0j ���   j j j j j Vj"�q�Ѓ�(^� �����������̋D$V�P�0� �R�@0j ���   j j j j j Vj5�q�Ѓ�(^� �����������̋D$V�P�0� �R�@0j ���   j j j �t$ j Vj<�q�Ѓ�(^� ���������̡ �V�@0j ���   j j j j �t$ ��j �t$$j�v�С ��t$8�@0�v�@t�Ѓ�0^� ��������̡ �j �@0j ���   j j j j j j j�q�Ѓ�(�������̡ �j �@0j ���   j j j j �t$j j�q�Ѓ�(� ��̡ �j �@0j ���   j j j j j j j�q�Ѓ�(�������̡ �j �@0j ���   j j j j j �t$ j�q�Ѓ�(� ��̡ �j �@0j ���   j j j j �t$ �t$ j&�q�Ѓ�(� ̡ �j �@0j ���   j j j j j j j(�q�Ѓ�(�������̡ �j �@0j ���   j j j j j j j#�q�Ѓ�(�������̡ �j �@0j ���   j j �t$�t$j �t$ j+�q�Ѓ�(� ��������������̡ �j �@0j ���   j j j j j j j0�q�Ѓ�(�������̡ ��t$�@0�q���   �Ѓ�� ���j�hNod�    P��V�P�3�P�D$d�    ���t$D�L$����� ��t$0�@h8kds�@4�L$�D$,    �С ��L$DQ�L$Qj �t$L�D$T    �t$L�@0�t$L���   �t$L�t$Hj2�v�Ћt$l��(�L$�D$$����薜���ƋL$d�    Y^�� � ̡ ��q�@0���   �Ѓ����������̋I��u3�� � �j �@0j ���   j j j j j �t$ j-Q�Ѓ�(� ��������̃�� �W�@j ���   ���L$(j�ЋL$$�D$� �j �@j���   �ЉD$� ��L$�@0Q�@`�L$Q�w�С ��T$�H0�D$,�pR�T$,R�T$$R�T$0R�0�Ah�w�Ѓ�(�|$( _t.�|$( t.�L$�T$;�~C�D$�;�}9�$�T$;�~.�D$��|$( u�L$�T$;�~�D$�;�}�   ��� 3���� ��SV�t$W��u�q� ��\$�@j ���   hdiuM���Ћ���tH;>u_^3�[� � �j �@hIicM���   ����;�u� �j �@h1icM���   ���Шu��>_^�   [� ������������j�hqod�    P��V�P�3�P�D$d�    � ��t$,�@hfnic�@T���ЋЅ�t� �j
�A�ʋ��   �Ѕ���   hfnic�D$P���(  �t$0P���D$(    �,����L$�D$$��������� ��΋@�@ �Ѓ��t� ��΋@�@ �Ѕ�u� �hfnic�@�΋@$�С ��t$4�@j
�@8���ЋL$d�    Y^�� ����������̡ ��q�@0���   �Ѓ�����������j�h�od�    P��$V�P�3�P�D$,d�    ��hmnrs�L$����� ��t$@�@j�@4�L$ �D$<    �ЍD$P�t$@�D$P������P� ��D$8���   �@8�Ћ ������   �D$�	P�D$< �у��L$�D$4�����ј���ƋL$,d�    Y^��0� ������������j�h�od�    P��$V�P�3�P�D$,d�    ��|$@ �SSSS�DSSSE�P�L$�.���� ��L$�@�D$4    �@ �Ћ �j�QP�B4�L$ �ЍD$P�t$@�D$P�������P� ��D$8���   �@8�Ћ ������   �D$�	P�D$< �у��L$�D$4���������ƋL$,d�    Y^��0� ���������������V��V��� �h�� �@0� �Ѓ��F�F    ���F   �F    ��^�V��N����t� �Q�@0�@�Ѓ��F    ^�������V��N�F    ��tk� �j �@0j ���   j j j j j j jQ�С ��t$<�H0�t$<3�9D$H�t$<���t$<j ��
P�v���   �Ѓ�D��t�~ t	�   ^� 3�^� �������������̋D$�A�I��u3�� � �Q�@0�@�Ѓ�� ��������̡ �S�@�\$�@ V�����=ckhc��   tz=cksata=TCAb��   � �W�@j ���   hdiem���Ћ��SW���F   �R�~ ��t��t��u3�������P�L���_^��[� �~ tg����P^[� �~ tU� �j �@0j ���   j j j j j j j �v�Ѓ�(��t)�F    ^�   [� =atnit�t$��S�\���^[� ^3�[� U��} ��   S�\$V�t$W�|$$��wy�$�|� 9t$��   �f9t$��   �Z9t$��   �N9t$��   �B�D$;�~:;���   �0�D$;�|(;�~~�"�D$;�|;�|p��D$;�~;�~b�9t$uZ� �j �@0j ���   j j j j j �t$0j�u��fn������(j���D$fn�����$S�Fm  ���E    _^[]� ��� �� �� ̡ ء � �� � � W��� �\  V�t$����   �$�� �D$f/D$�4  ��   �D$f/D$�  ��   �L$f/L$�  �   �L$f/L$��   �   �T$f/T$��   �D$$f/���   �n�T$f/T$r`�D$$f/���   �N�T$f/T$r@�D$$f/���   �.�T$f/T$v �D$$f/�sl��D$f.D$���DzX� �j �@0j ���   j j j j j �t$(j�w���D$L��(�t$,���D$�D$0�$V�k  ���G    ^_�$ �I ¢ ٢ � � � B� b� �� �� �������������D$j���D$�D$0�D$�D$(�$�t$$�t$$�+����  ���������D$j���D$�D$0�D$�D$(�$�t$$�t$$������  ���������D$j���D$�D$0�D$�D$(�$�t$$�t$$�����  ��������V��V��� �h�� �@0� �Ѓ��F�F    �<��F   ��^��������V��N����t� �Q�@0�@�Ѓ��F    ^������̡ �V�@��L$�@ ��=cksat]=ckhct�t$���t$�/���^� j j j j j j �F   � �j �@0j ���   j �v�Ѓ�(��t!�F    �   ^� �~ t����P^� 3�^� �j�h�od�    PQV�P�3�P�D$d�    ��t$��� �V�@0h�� � �Ѓ��F�F    �F   �D$ �L$�d��F� �j �@hmyal���   �D$    �ЉF��t��t�F    � ��L$�@j
���   hhfed�ЉF�ƋL$d�    Y^��� ����̡ �V�@��L$�@ ��=ytsdt�t$���t$�v���^� � ��v�@0���   �Ћ�����P�   ^� ������������3���������������3�������������������������������3���������������3���������������3���������������3�� �����������Q�L$�$    ��n���D$Y� ������̋A��uË ���������������������V���PD��t�D$9Ft
�F����PH^� ������������̋A�������������j0�t$�a  ����j0�t$��z����P�la  �����������j�hpd�    P���P�3�P�D$d�    �t$(�D$�t$(P�z��j0P�D$0    �a  � ��L$�@Q�@�D$4�����Ѓ��L$d�    Y�����������������j�h0pd�    P���P�3�P�D$d�    �t$,�D$�t$,�t$,P��{��j0P�D$4    �`  � ��L$�@Q�@�D$8�����Ѓ��L$d�    Y�������������j$�t$�U`  3Ƀ���������������j$�t$�y����P�,`  3Ƀ����������������������j�hSpd�    P��S�P�3�P�D$d�    �t$,�D$�t$,P�Zy��j$P�D$4    ��_  � �3ۋI���I�D$P���D$8�����у��ËL$d�    Y[����j�hvpd�    P��S�P�3�P�D$d�    �t$0�D$�t$0�t$0P�z��j$P�D$8    �F_  � �3ۋI���I�D$ P���D$<�����у��ËL$d�    Y[���������������̡ ��t$�@�t$���   j �Ѓ�����t$� ��t$�@�t$���   j �Ѓ���������������̡ ��@���  �� ��@0���   ��j�h�pd�    P��VW�P�3�P�D$ d�    �t$8�D$    � ��t$8�@0�L$���   Q�Ћ�� ��|$<�IW�I�D$8   �ѡ �W�@V�@�Ћ ��D$(�IP�I�D$(   �D$D �у��ǋL$ d�    Y_^�� ����j�h�pd�    P��(SUVW�P�3�P�D$<d�    �D$    � ��|$L�@W�@�D$H    �Ѓ�� ��L$P�@3ۋ��   SS�D$L    �D$    �ЋL$P�D$� �S�@j���   �Ћ����&  3���I ��~|� ��L$�@Q�@�С �j �@j��@�L$(h��Q�Ѓ�� ��ϋ@�D$D   �@<�Ћȡ �j��@j��@L�T$$RQ���С ��L$�@Q�@�D$H �Ѓ�V�t$�D$4P�!������� ��ϋ@�D$D   �@<�Ћȡ �j��@j��@LVQ���С ��L$,�@Q�@�D$H �С ��L$T�@�����   j ��
UC�ЉD$� �j �P�M���   Q�L$X�ҋ���������ǋL$<d�    Y_^][��4�����������̡ ��@0���   �� ��@0���   �� ��@0���   ����W��JR��A(�P$j j h����_  �������������̸�������������j�hAqd�    P��8SVW�P�3�P�D$Hd�    ����L$Q���P(���W�D$P    ��t&� �j �A0j ���   j j j j Vj jR�Ѓ�(� ��L$�@Q�@�D$T�����С ��L$�@Q�@�Ѓ��O�D$P   ��t'� �j �@0j ���   j �T$ Rj jj?j Q�Ѓ�$� ��L$�@Q�@�D$T�����С ��L$�@Q�@�Ѓ��O�D$P   ��u3��>� ��T$Rj j j h  
 j�T$,R�D$,    �@0h�  ���   jQ�ЋD$8��(��� ��L$�@Q�@���D$T�����Ѓ���t3��L$Hd�    Y_^[��Dá ��L$�@Q�@�Ѓ��O�D$P   ��t'� �j �@0j ���   j �T$ Rj j j8j Q�Ѓ�$� ��L$�@Q�@�D$T�����ЋO����t� �j�@0Q�@P�Ѓ��L$4�z������ ��D$$�IP�I�D$T   �у�Vh   h  K j;�D$4Ph	��h�  ���D$l�R���� ��L$$�@Q�@�D$T�Ѓ��L$4�D$P�����g����O��t� �Q�@0�@X�Ѓ��O��t� �Q�@0�@X�Ѓ��O��t&� �j �@0j ���   j j j jj j jQ�Ѓ�(j�$��W  ���   �L$Hd�    Y_^[��D������j�hdqd�    P��VW�P�3�P�D$$d�    ��j�N��v  �F4    �F8    �F<    W��F(� �h�   �@0�v�@�С ��L$�@Q�@�С �j �@j��@�L$(h��Q�Ѓ�j j �D$P�D$P���D$<    �D$�  �D$     谿��� ��L$�@Q�@�D$0�����Ѓ��Nj j��u  �L$$d�    Y_^��$������j�h�qd�    P��\VW�P�3�P�D$hd�    �� ��L$�@Q�@�С �j �@j��@�L$ h�Q���F(�YȖǄ$�       �D$ �  �D$$    �,�P�D$LP�E  �L$0QP�D$HPƄ$�   ��  ��(j j P�D$P��Ƅ$�   豾��� ��L$$�@Q�@�D$t�С ��L$8�@Q�@�D$x �С ��L$�@Q�@�D$|�����Ѓ��L$Thtats舃��� �j�@j�@0�L$\�D$x   �С ��F(�@�@,���L$\�$j�ЍD$TP�D$P�D$LP���D$�  �D$    ����� ��L$D���   Q� �Ѓ��~4 t_� ��N0�@P�@h�ЋF4��t�v8�Ѓ��F<�F8    �F4    �� �h��@h�  ��0  �Ѓ�� ��N0�@P�@l�ЍL$T�D$p�����؂���L$hd�    Y_^��h� ����j�h�qd�    P��@VW�P�3�P�D$Ld�    �� ��|$\�@�ϋ@ ��=MicM��   =ckhctg=fnic�9  j�L$<�����L$`P�D$X    �\����L$8�D$T�����;���� ��L$`�@j�@4j�и   �L$Ld�    Y_^��L� ����P����؋L$Ld�    Y_^��L� � �j �@hIicM���   ����=�����   htats�L$(�z���� �j �@j�@0�L$,�D$\   �ЍD$$P�D$P�D$P���D$�  �D$    ����� ��L$���   Q� �Ѓ��L$$�D$T�����O����N�F   ��t� �Q�@0�@�Ѓ��t$`��W�����L$Ld�    Y_^��L� �l$V��t3�^� j�N�&r  j��R  �N���F    ��t� �Q�@0�@�Ѓ��   ^� ����j����q  j�R  ��3������������D$�A(� �̍A�������������VW��~4 tC��    � �h���@h~  ��0  ��j
�/]  � ��v �@P�@�Ѓ���uM9F4uá ��N0�@P�@h�Ѓ~4 t9� �hȔ�@h�  ��0  �С ����@P�N0�@l���o���_3�^� �D$�F8�D$�F4� �S�@P�N0�@l�Ѓ~4 t#j
�\  � ��v �@P�@�Ѓ���u89F4uݡ ��N0�@P�@h�Ћ~<�F<    � ��N0�RP�Rl��[��_^� [_3�^� �j�h�qd�    P��V�P�3�P�D$d�    �L$��~���L$0� ��D$$    ��t"�@4Q�@�Ѓ���t'��L$Q�t$8���R(�'�@0�t$,�@�Ћȃ���u3��?��T$R�t$8�P �� ��L$�@�@ �Ѓ��t� ��L$�@0Q�t$0�@x�Ѓ��L$�D$$�����~���ƋL$d�    Y^�� á �V�@j �t$���   ��L$�Ћ���u�    �F^� ��u9Ft�   ^� ������������V�t$W��;t$u� ��L$�@j ���   htsem�Ѕ�u`� ��L$�@j ���   hrdem�Ѕ�uA�D$�D$�H��t2� �j �@0�T$�@,RVQ�Ѓ���t�t$���	  _�   ^� _3�^� ������������j�h rd�    P��0VW�P�3�P�D$<d�    ��� ��L$�@Q�@�С ��L$ �@Q�@�D$L    �Ѓ��L$L�D$P�t$T�D$4P�D$P�~z���Ћ ��D$D�A�L$�@QR�С ��L$4�@Q�@�D$P�С ��L$(�@Q�@�D$T �С ���@V�@�С ��L$ �@V�@Q�Ѓ�����	  � ��L$�@Q�@�D$H�����Ѓ��L$<d�    Y_^��<� �������j�hCrd�    P��SV�P�3�P�D$$d�    �ًt$<;t$@��   � ��L$8�@j ���   htsem�Ѕ���   � ��L$8�@j ���   hrdem�Ѕ���   � ��L$�@Q�@�Ѓ��L$4�D$P�D$P�D$4    �t$�D$    虹����u3��5� ����@��@V�С ��L$(�@V�@Q�Ѓ����  �   � ��D$�IP�I�D$0�����у��ƋL$$d�    Y^[��$� 3��L$$d�    Y^[��$� �̡ �V�@j �t$���   ��L$�Ћ���u�    �F^� ��u9Ft�   ^� �����������̃�V�t$W��;t$ uy� ��L$�@j ���   htsem�Ѕ�uZ� ��L$�@j ���   hrdem�Ѕ�u;�L$�D$�D$�D$P�D$P�t$������t�t$���S  _�   ^��� _3�^��� �����������̃�� �V�@�����   W��$�t$��L$���\$����u�D$�    �F^��� ��u�Ff.D$���D{�   ^��� �̃�SV�t$��;t$ ��   � ��L$�@j ���   htsem�Ѕ�ur� ��L$�@j ���   hrdem�Ѕ�uS�D$W��H�D$��t?� �j �@0�T$�@0RVQ�Ѓ���t"�D$�����$�W  ^�   [��� ^3�[��� ��0� �V��W��L$Q�t$@�D$�D$�D$�@�L$$���   Q�L$D���~�~P�~H����uf�^f�V�    f�N^��0� ��u3�Ff.ß��Dz�Ff.��Dz�Ff.����D{�   ^��0� ���̃�4�D$@S�\$HV�t$TW�|$T�L$;�t;�t;���   � ��L$H�@j ���   htsem�Ѕ���   � ��L$H�@j ���   hrdem�Ѕ���   �L$D�D$�D$�D$$�D$(P�D$P�D$ PW��D$,P�D$8�D$@�D$H�t$ �|$(�\$0�������t<�~D$(�L$����f� �~D$Hf�@�~D$Pf�@��  �   _^[��4� _^3�[��4� ����������̃�0� �V��W��D$����L$Q�t$@�D$�@�L$,���   Q�L$D���~ �~H�f�D$f�L$���uf�F�    f�N^��0� ��u�D$P�FP��   ����t�   ^��0� �������̃�SV�t$0��;t$4��   � ��L$(�@j ���   htsem�Ѕ���   � ��L$(�@j ���   hrdem�Ѕ�uh�L$$�D$�D$P�t$0W��D$����D$P�D$$�t$������t.�~D$���ċ�f� �~D$(f�@��  �   ^[��� ^3�[��� ������̃�V�t$W�|$ �f.���Dz�Ff.G���D{a�G�Y����D$�D$�$藟  �F�\$�Y�D$�D$�$�x�  �D$�\$��f.D$���D{_�   ^���_3�^���������������j�hyrd�    PQV�P�3�P�D$d�    �D$    � ��t$�@V�@�D$    �С �V�@�t$(�@�Ѓ�� ��΋@�D$    �@<�D$   �Ћ �j��Qj��t$,�RLP���ҋƋL$d�    Y^���������������V��N����t� �Q�@0�@�Ѓ��D$�F    t	V�{\������^� ��V��~ ���u� ��v�@4� �Ѓ��D$�F    �F    t	V�4\������^� ����������̋���u�D$�    �A� ��u�A;D$t�   � ��̋���u�D$�    �A� ��u�Af.D$���D{�   � ������̋���u*�~D$f�A�~D$f�A�~D$�    f�A� ��u9�Af.D$���Dz"�Af.D$���Dz�Af.D$���D{�   � ���������������V�����u �~D$f�F�~D$�    f�F^� ��u�D$P�FP���������t�   ^� ���j�h�rd�    PV�P�3�P�D$d�    ���D$    ���u!�    � ��N�@Q�@�L$Q�Ѓ��#��u� ��T$�@�N�@xR�Ѕ�t�   � ��L$�@Q�@�D$�����Ѓ��L$d�    Y^��� ����������j�h�rd�    P���P�3�P�D$d�    �t$0�D$    � ��T$�@R�@P�ЋL$,P�D$(   �q���L$�D$   �D$$ �q���D$,�L$d�    Y��$� �j�h1sd�    P�� �P�3�P�D$$d�    �t$<�D$    � ��t$<�@�T$���   R�ЋL$4P�D$0   ��  �L$�D$   �D$, �`  �D$4�L$$d�    Y��,� ����������j�h�jd�    P��VW�P�3�P�D$ d�    �t$4�D$    � ��L$�@Q�@(�Ћ�� ��|$8�IW�I�D$4   �ѡ �W�@V�@�Ћ ��D$$�IP�I�D$$   �D$@ �у��ǋL$ d�    Y_^�� ����������̋L$�D$Q��D$j�t$�A�L  �����������������̸   �����������V�t$��t���u7j�t$��K  ����u3�^Ë��K  �ȅ�t��t��D$3�;AOʋ�^���������Vj j�t$����������t�@��t����^� 3�^� ����Vj j�t$���p�������t�@��t����^� 3�^� ����Vj j�t$���@�������t�@��t����^� ����������Vj j�t$����������t�@��t����^� 3�^� ����Vj j�t$�����������t�@��t����^� 3�^� ����Vj j�t$����������t�@��t����^� 3�^� ����Vj j �t$����������t�@ ��t�t$����^� 3�^� j�hysd�    P��4VW�P�3�P�D$@d�    ��j j$�t$\�D$    �$�������to�@$��th�L$(Q���Ћ���|$Pj ��W�D$L   �    �B    � ����   �FP�AR�Ћ ��D$<���   P�	�D$   �D$X �ы��g�L$�EM���t$P�D$��Nj �    �A    � ��T$���   R�@Q�D$T   �Ћ ��D$$���   P�	�D$   �D$X �ыƃ��L$@d�    Y_^��@� Vj j(�t$��� �������t�@(��t�t$����^� ������Vj j,�t$�����������t�@,��t����^� 3�^� ����Vj j0�t$�����������t�@0��t����^� 3�^� ���̋D$�@�< �@�� �@�� �@�< �@�� �@�� �@ �� �@$�< �@(�� �@,�� �@0�� �@4�� ��������3�� ��`T��`$��`0��`4��`8��`<��`D��`L��`P�������������̋D$� �� ��������������������̡ ��@$�@X����̡ ��@$�@\������t$� ��t$�@$�t$�@`Q�Ѓ�� j�h�sd�    PQV�P�3�P�D$d�    ��t$� �V�@�@�С �V�@$�D$    �@D�Ѓ��ƋL$d�    Y^�����������������j�h�sd�    PQV�P�3�P�D$d�    ��t$� �V�@�@�С �V�@$�D$    �@D�С ��t$$�@$V�@d�Ѓ��ƋL$d�    Y^��� ����������j�h�sd�    PQV�P�3�P�D$d�    ��t$� �V�@�@�С �V�@$�D$    �@D�С ��t$$�@$V�@�Ѓ��ƋL$d�    Y^��� ����������j�htd�    PQV�P�3�P�D$d�    ��t$� �V�@�@�С �V�@$�D$    �@D�С �V�@$�t$(�@L�Ѓ��ƋL$d�    Y^��� ����������j�h4td�    PQV�P�3�P�D$d�    ��t$� �V�@$�D$    �@H�С �V�@�D$�����@�Ѓ��L$d�    Y^����������̡ ��t$�@$Q�@L�Ѓ�� �������̡ ��@$�@����̡ �Q�@$�@�Ѓ����������������j�hptd�    P��VW�P�3�P�D$ d�    �D$    � �Q�@$�L$�@Q�Ћ�� ��|$8�IW�I�D$4   �ѡ �W�@V�@�Ћ ��D$$�IP�I�D$$   �D$@ �у��ǋL$ d�    Y_^�� � ����������̡ ��t$�@$Q�@�Ѓ�� ��������j�h�td�    P�� VW�P�3�P�D$,d�    �D$    � �Q�@$�L$�@ Q�Ћ�� ��|$D�IW�I�D$@   �ѡ �W�@$�D$D�@D�С �W�@$V�@L���D$$   � ��L$(�@$Q�@H�D$P   �Ћ ��D$,�IP�I�D$T �у� �ǋL$,d�    Y_^��,� ��������������j�hud�    P�� VW�P�3�P�D$,d�    �D$    � �Q�@$�L$�@$Q�Ћ�� ��|$D�IW�I�D$@   �ѡ �W�@$�D$D�@D�С �W�@$V�@L���D$$   � ��L$(�@$Q�@H�D$P   �Ћ ��D$,�IP�I�D$T �у� �ǋL$,d�    Y_^��,� ��������������j�hLud�    P�� �P�3�P�D$$d�    �D$P�D$    ������t$4���D$0   �(����D$   � ��L$�@$Q�@H�D$0   �Ћ ��D$�IP�I�D$4 �ыD$<���L$$d�    Y��,� ����̡ �Q�@$�@(��Yá �Q�@$�@h��Yá ��t$�@$Q�@,�Ѓ�� �������̡ ��t$�@$Q�@0�Ѓ�� �������̡ ��t$�@$Q�@4�Ѓ�� �������̡ ��t$�@$Q�@8�Ѓ�� �������̡ ��t$�@$�t$�@PQ�Ѓ�� ���̡ ��t$�@$Q�@T�Ѓ�� �������̡ ��@$�@l����̡ ��@$�@p����̡ �V�@$��@LV�t$�Ѓ���^� ��j�h�ud�    PQV�P�3�P�D$d�    �D$    � ��t$�@V�@�D$    �С �V�@$�D$   �@D�С �V�@$�t$,�@L�Ћ ��t$4�I$V�I@�D$,    �D$    �у��ƋL$d�    Y^�������������̡ �V�@$�t$�@@��V�Ѓ���^� �̡ ��t$�@$Q�@<�Ѓ�� �������̡ ��t$�@$Q�@<�Ѓ����@� ���j�h�ud�    P��VW�P�3�P�D$ d�    �D$    � �Q�@$�L$�@tQ�Ћ�� ��|$8�IW�I�D$4   �ѡ �W�@V�@�Ћ ��D$$�IP�I�D$$   �D$@ �у��ǋL$ d�    Y_^�� � ����������̡ ��@(�@����̡ ��@(�@����̡ ��@(�@����̡ ��@(�@����̡ ��@(�@ ����̡ �j�t$�@(�t$�@��� �������t$� ��t$�@(�t$�@$��� ���̡ ��@(�@(����̡ ��@(�@,����̡ ��@(�@0����̡ ��@(�@4����̡ ��@(�@X����̡ ��@(�@\����̡ ��@(�@`����̡ ��@(�@d����̡ ��@(�@h����̡ ��@(�@l����̡ ��@(�@p����̡ ��@(�@t����̡ ��@(�@x����̡ ��@(���   ��j�h�ud�    P��V�P�3�P�D$d�    �� ��L$�@Q�@�Ѓ��D$P���D$$    �   ��u3��� ��L$�@$Q�t$,�@�Ѓ��   � ��D$�IP�I�D$$�����у��ƋL$d�    Y^��� ��������Q� ��T$�@(R�@X�Ѕ�uY� �D$3�8L$����   Y� �������������j�h
vd�    P��V�P�3�P�D$ d�    �� ��D$    �D$    �@(�L$�@hQ���Ѕ���   �L$� ���uM�@�L$�@Q�С ��t$4�@�L$�@Q�D$4    �С ��L$�@Q�@�D$8�����Ѓ��   �@h����   hj  Q�Ћȡ ����L$�@(��u�@4j�����3��L$ d�    Y^��$� �@j �t$Q���Ѕ�u"�D$P�H����3��L$ d�    Y^��$� � �j �H�D$HP�t$�A�t$<�ЍD$P��G�����   �L$ d�    Y^��$� ����̡ �V�@(W�|$�@pW���Ѕ�t8� ��΋P(�GP�Bp�Ѕ�t!� ��΋P(�GP�Bp�Ѕ�t
_�   ^� _3�^� ������̡ �V�@(W�|$�@tW���Ѕ�t8� ��΋P(�GP�Bt�Ѕ�t!� ��΋P(�GP�Bt�Ѕ�t
_�   ^� _3�^� ������̡ �S�@(V�@pW�|$W���Ѕ���   � ��΋P(�GP�Bp�Ѕ���   � ��΋P(�GP�Bp�Ѕ�tn� ��_�@(S�@p���Ѕ�tW� ��΋P(�CP�Bp�Ѕ�t@� ��΋P(�CP�Bp�Ѕ�t)�GP��������t�G$P��������t_^�   [� _^3�[� ��������̡ �S�@(V�@tW�|$W���Ѕ���   � ��΋P(�GP�Bt�Ѕ���   � ��΋P(�GP�Bt�Ѕ�tn� ��_�@(S�@t���Ѕ�tW� ��΋P(�CP�Bt�Ѕ�t@� ��΋P(�CP�Bt�Ѕ�t)�G0P���/�����t�GHP��� �����t_^�   [� _^3�[� ��������̡ ��@(�@8����̡ ��@(�@<����̡ ��@(�@@����̡ ��@(�@D����̡ ��@(�@H����̡ ��@(�@L����̡ ��D$�@(Q�@P�$��� ���̡ ��D$�@(���@T�$��� �̡ ��t$�@(�t$�@|��� �������̡ ��t$�@(�t$���   ��� �����j�h-vd�    P��V�P�3�P�D$d�    ��L$(�D$P����P���D$$    �\   � ����I�D$�IP�D$$�����у��ƋL$d�    Y^��� ������̡ ��|$ �P(�����D$�B8������Q� �V�@W�@d���L$j �Ћ �h��I�p���   h�  V�ыȡ ����L$��u�@(j��@4����_3�^Y� �@j �@hVQ�L$�С �V�@(�ϋ@H�Ѕ�t2� �V�@(�t$�@ ���Ѕ�t�D$P�   �8C������_^Y� �D$P3��!C������_^Y� �����̡ �V�@(W�|$�@P�Q���$�Ѕ�tF� ��G�@(Q�@P���$�Ѕ�t(� ��G�@(Q�@P���$�Ѕ�t
_�   ^� _3�^� � �V�@(W�|$�@T������$�Ѕ�tJ� ��G�@(���@T���$�Ѕ�t*� ��G�@(���@T���$�Ѕ�t
_�   ^� _3�^� ���������̡ �V�@(W�|$�@P�Q���$�Ѕ��  � ��G�@(Q�@P���$�Ѕ���   � ��G�@(Q�@P���$�Ѕ���   � ��G�@(Q�@P���$�Ѕ���   � ��G�@(Q�@P���$�Ѕ���   � ��G�@(Q�@P���$�Ѕ�ts� ��G�@(Q�@P���$�Ѕ�tU� ��G�@(Q�@P���$�Ѕ�t7� ��G �@(Q�@P���$�Ѕ�t�G$P���������t
_�   ^� _3�^� ��������̡ �V�@(W�|$�@T������$�Ѕ���   � ��G�@(���@T���$�Ѕ���   � ��G�@(���@T���$�Ѕ���   � ��G�@(���@T���$�Ѕ�th� ��G �@(���@T���$�Ѕ�tH� ��G(�@(���@T���$�Ѕ�t(�G0P���T�����t�GHP���E�����t
_�   ^� _3�^� � ��@(� �����̡ �V�@(�t$�@�6�Ѓ��    ^�̡ ��@(���   �� ��@(�@����̡ ��@(�@����̡ �V�@(�t$�@�6�Ѓ��    ^�̡ ��t$�@,�t$�@Q�Ѓ�� ���̡ ��@,�@����̡ ��@,�@����̡ ��@,�@����̡ ��@,�@ ����̡ ��@,�@(����̡ ��@,�@$����̡ ��@,�@�����j�hyvd�    P�� VW�P�3�P�D$,d�    �D$    � ��T$�@,R�@�Ћ�� ��|$<�IW�I�D$8   �ѡ �W�@$�D$<�@D�С �W�@$V�@L���D$   � ��L$ �@$Q�@H�D$H   �Ћ ��D$$�IP�I�D$L �у��ǋL$,d�    Y_^��,� ��������������̡ �j �@,j � �Ѓ�������������̡ �V�@,�t$�@�6�Ѓ��    ^�̡ ��@,�@4����̡ ��@,�@8�����j�h�vd�    P�� VW�P�3�P�D$,d�    �D$    � ��T$�@,R�@<�Ћ�� ��|$<�IW�I�D$8   �ѡ �W�@$�D$<�@D�С �W�@$V�@L���D$   � ��L$ �@$Q�@H�D$H   �Ћ ��D$$�IP�I�D$L �у��ǋL$,d�    Y_^��,� ���������������j�hwd�    P��VW�P�3�P�D$ d�    �t$4�D$    � ��T$�@,R�@@�Ћ�� ��|$0�IW�I�D$,   �ѡ �W�@V�@�Ћ ��D$�IP�I�D$   �D$8 �у��ǋL$ d�    Y_^�� � �������̡ ��@,�@,����̡ �V�@,�t$�@0�6�Ѓ��    ^�̡ ��@���  �� ��@���  �� ��@���  �� ��@���  �� ��@�@����̡ ��@�@����̡ ��@�@����̡ ��@�@����̡ ��@�@����̡ ��@�@����̡ ��t$�@�t$�@\��� �������̡ ��t$�@�t$��  ��� ����̡ ��D$�@���@ �$��� �̡ ��D$�@Q�@$�$��� ���̡ ��D$�@���@(�$��� �̡ ��@�@,����̡ ��@�@0����̡ ��@�@4����̡ ��@�@8����̡ ��@�@<����̡ ��@�@@����̡ ��@�@D����̡ ��@�@H����̡ ��@�@L����̡ ��@�@P����̡ ��@���   �� ��t$�@Q��  �Ѓ�� ����̡ ��@�@T����̡ ��@�@X����̋T$��u3�� � �R�@ Q�@(�Ѓ��   � ��������̡ ��@���   �� ��@�@`����̡ ��@�@d����̡ ��@�@h����̡ ��@�@l����̡ ��@�@p����̡ ��@�@t����̡ ��@���   �� ��@��  �� ��@�@x����̡ ��@�@|����̡ ��@���   �� ��@���   �� ��@���   �� ��@���   �� ��@���   �� ��@���   �� ��@���   �� ��@���   �� ��@���   �� ��@���   �� ��@���   �� ��@���   �� ��t$�@Q��  �Ѓ�� ����̡ ��@���   �� ��@���   ���T$��t� �R�@ Q�@$�Ѓ���t�   � 3�� ����̡ �Q�@ �t$�@L�t$�Ѓ�� ���̡ ��@���   �� ��@���   �� ��@���   �� ��@���   �� ��@���   �� ��@���   �� ��@���   �� ��@���   �� ��@���   �� ��@���   �� ��@���   �� ��@���   �� ��@���   �� �V�@�t$���   V�Ѓ��    ^���������������̡ ��@� �����̡ ��@�@����̡ ��@���   �� ��@��   �� ��@�@����̡ ��@�@����̡ ��@�@����̡ ��@�@����̡ ��@�@����̡ ��@���  �� ��@�@�����j�h,wd�    P��V�P�3�P�D$$d�    �t$4�D$P������� ��L$�@$Q�@�D$0    �Ѓ���t_� ��L$�@j�@Q�Ѓ���u�D$P��������t3� �j�@V�@�Ѓ���u� �V�@�@�Ѓ���t�   �3�� ��L$�@$Q�@H�D$0   �Ћ ��D$�IP�I�D$4�����у��ƋL$$d�    Y^��(���������������̡ ��@�@ ����̡ ��@�@(����̡ ��@��  �� ��@��   �� ��@��  �� ��@��  ��j�hxwd�    P�� VW�P�3�P�D$,d�    �D$    � ��L$�@Q�@$�Ћ�� ��|$@�IW�I�D$<   �ѡ �W�@$�D$@�@D�С �W�@$V�@L���D$    � ��L$$�@$Q�@H�D$L   �Ћ ��D$(�IP�I�D$P �у��ǋL$,d�    Y_^��,��j�h�wd�    P�� VW�P�3�P�D$,d�    �D$    � ��L$�@Q���  �Ћ�� ��|$@�IW�I�D$<   �ѡ �W�@$�D$@�@D�С �W�@$V�@L���D$    � ��L$$�@$Q�@H�D$L   �Ћ ��D$(�IP�I�D$P �у��ǋL$,d�    Y_^��,���������������Qj�t$�D$    �  �D$�������j�hJxd�    P��<SVW�P�3�P�D$Ld�    �D$    �H���t�D$0P�^������D$T   �   �@� ��L$�@Q�@�С ��L$�@$Q�@D�D$\   �Ѓ��|$�D$T   �   � ��t$\�@V�@�\$�С �V�@$�D$\   �@D�С �V�@$W�@L�Ѓ�����t;����\$� ��L$�@$Q�@H�D$X   �С ��L$�@Q�@�D$\�Ѓ��D$T    ��t<����\$� ��L$0�@$Q�@H�D$X   �Ћ ��D$4�IP�I�D$\ �у��ƋL$Ld�    Y_^[��H���������������j�h�xd�    P�� VW�P�3�P�D$,d�    �t$@�D$    � ��L$�@Q���  �Ћ�� ��|$D�IW�I�D$@   �ѡ �W�@$�D$D�@D�С �W�@$V�@L���D$$   � ��L$(�@$Q�@H�D$P   �Ћ ��D$,�IP�I�D$T �у� �ǋL$,d�    Y_^��,����������̡ ��@��D  �� ��@��H  �� ��@��L  ��j�h�xd�    P��VW�P�3�P�D$ d�    �t$8�D$    � ��t$8�@�L$���  Q�Ћ�� ��|$<�IW�I�D$8   �ѡ �W�@V�@�Ћ ��D$(�IP�I�D$(   �D$D �у��ǋL$ d�    Y_^�� ���̡ ��@���  �� ��@���  �� �Q���   �@X�Ћȃ���u� � ��t$�@|�t$�@Q�Ѓ�� ������̡ �Q���   �@X�Ћȃ���u� � ��t$�@|�t$�@8Q�Ѓ�� ������̋T$V��j �� �j �@j �@R�Ѓ��F��^� ������̡ �V�@j �@j ��j �6�Ѓ��F^�V��N��u3�^� � �Q�t$�@�t$�@�6�Ѓ��F�   ^� ��������̋D$V�0W�9;�t_3�^� �P��u��u9pu9qu��u�9yu�_�B^� S�Y��u!��u9yu��u2��u.9pu)[_�   ^� ��t��t;�u�P��t�A��t�;�t�[_3�^� �������t$�g������@� ���������������Vh(�j\hD ����������t�@\��tV�Ѓ���^�����Vh(�j\hD ���\�������t3�@\��t,V��h(�jxhD �:�������t�@x��t
V�t$�Ѓ���^� �����������̃�Vh(�j\hD �����������tL�@\��tEV�ЋD$h(�jdhD �D$�D$    �D$    ��������t�@d��t�L$QV�Ѓ���^��� �������������Vh(�j\hD ���|�������t3�@\��t,V��h(�jdhD �Z�������t�@d��t
�t$V�Ѓ���^� ������������Vh(�j\hD ����������t\�@\��tUV��h(�jdhD ���������t�@d��t
�t$V�Ѓ�h(�jhhD ���������t�@h��t
�t$V�Ѓ���^� ���Vh(�j\hD ������������   �@\��t~V��h(�jdhD �v�������t�@d��t
�t$V�Ѓ�h(�jhhD �M�������t�@h��t
�t$V�Ѓ�h(�jhhD �$�������t�@h��t
�t$V�Ѓ���^� ������Vh(�j`hD �����������t�@`��tV�Ѓ�^�������Vh(�jdhD ����������t�@d��t
�t$V�Ѓ�^� Vh(�jhhD ����������t�@h��t
�t$V�Ѓ�^� Vh(�jlhD ���\�������t�@l��tV�Ѓ�^�������Vh(�jphD ���,�������t�@p��t�t$V�Ѓ�^� �,�^� �������Vh(�jxhD �����������t�@x��t
V�t$�Ѓ���^� ��������������Vh(�j|hD ����������t�@|��tV�t$�Ѓ�^� 3�^� ����������Vh(�j|hD ���l�������t�@|��tV�t$�Ѓ����@^� �   ^� ��j�hyd�    P��V�P�3�P�D$d�    ��h(�jthD �D$    ��������tu�@t��tn�t$(�L$VQ�Ѓ��t$$P���D$    �`���h(�j`hD �D$   �D$( ��������tv�H`��to�D$P�у��ƋL$d�    Y^��� h(�j\hD �t����t$0����t4�@\��t-V��h(�jdhD �N�������t�@d��th,�V�Ѓ��ƋL$d�    Y^��� Vh(�h�   hD ���	�������t���   ��t�t$V�Ѓ�^� 3�^� ����Vh(�h�   hD �����������t���   ��t�t$V�Ѓ�^� 3�^� ����VW��3����$    �h(�jphD ��������t�@p��t	VW�Ѓ���,��8 tF��_��^�������SU�l$V��3�W�d$ h(�jphD �/�������t�@p��t	VS�Ѓ���,��8 tnh(�jphD ���������t�@p��tVU�Ѓ�����,�h(�jphD ���������t�@p��t	VS�Ѓ���,�W���Z�����tF�`����D$_��t�0��~=h(�jphD ��������t�@p��t	VS�Ѓ���,��8 u^]�   [� ^]3�[� �����������̃�Vh(�h�   hD ���&�������t?���   ��t5�t$�L$VQ��h(�j`hD ���������t�@`��t
�L$Q�Ѓ���^��� �������j�hMyd�    P��V�P�3�P�D$d�    h(�h�   hD �D$    ��������ty���   ��to�t$,�L$�t$,Q�Ѓ��t$$P���D$    �����h(�j`hD �D$   �D$( �;�������ts�H`��tl�D$P�у��ƋL$d�    Y^���h(�j\hD ������t$0����t3�@\��t,V��h(�jxhD ���������t�@x��t
V�t$,�Ѓ��ƋL$d�    Y^����������������̋���������������h(�jhD ��������t	�@��t��3��������������V�t$�> t+h(�jhD �E�������t�@��tV�Ѓ��    ^���������̃|$ W��t1h(�jhD ��������t�@��t�t$�t$W�Ѓ�_� 3�_� ���������������Vh(�jhD ����������t�@��t�t$V�Ѓ�^� 3�^� ����������Vh(�jhD ���|�������t�@��t�t$V�Ѓ�^� 3�^� ����������Vh(�j hD ���<�������t�@ ��tV�Ѓ�^�3�^���Vh(�j$hD ����������t�@$��tV�Ѓ�^�3�^���Vh(�j(hD �����������t�@(��t�t$�t$�t$V�Ѓ�^� 3�^� ��Vh(�j,hD ����������t�@,��t�t$�t$V�Ѓ�^� 3�^� ������Vh(�j(hD ���\�������t�@0��t�t$�t$�t$V�Ѓ�^� 3�^� ��Vh(�j4hD ����������t�@4��tV�Ѓ�^�3�^���Vh(�j8hD �����������t!�@8��t�t$�t$�t$�t$V�Ѓ�^� 3�^� ��������������Vh(�j<hD ����������t�@<��t
�t$V�Ѓ�^� Vh(�h�   hD ���i�������u^� �t$���   V�Ѓ�^� ����������Vh(�h�   hD ���)�������u^� �t$���   V�Ѓ�^� ����������Vh(�h�   hD �����������u^� �t$���   V�Ѓ�^� ����������Vh(�h�   hD ����������t�t$���   �t$�t$V�Ѓ�^� ������Vh(�jDhD ���l�������t�@D��tV�Ѓ�^�3�^���Vh(�jHhD ���<�������t�t$�@HV�Ѓ�^� ����Vh(�jLhD ����������u^� �t$�@LV�Ѓ�^� Vh(�jPhD �����������u^� �t$�@P�t$V�Ѓ�^� ������������Vh(�h�   hD ����������u^� �t$���   �t$�t$V�Ѓ�^� ��Vh(�h�   hD ���Y�������u^� �t$���   �t$�t$�t$�t$V�Ѓ�^� ����������Vh(�jThD ����������u^Ë@TV�Ѓ�^���������Vh(�jXhD �����������t�t$�@XV�Ѓ�^� ����j�h�yd�    P��V�P�3�P�D$ d�    ��h(�h�   hD �D$    �~�������t~���   ��tt�t$4�L$Q���Ћt$0P���D$,   �����h(�j`hD �D$   �D$4 �.���������   �H`����   �D$P�у��ƋL$ d�    Y^��$� h(�j\hD �D$     �D$$    �D$(    ������t$<����t4�@\��t-V��h(�jdhD ��������t�@d��t�L$QV�Ѓ��ƋL$ d�    Y^��$� ������������Vh(�h�   hD ���Y�������t���   ��t�t$���t$�t$��^� 3�^� ��������������Vh(�h�   hD ���	�������t���   ��t�t$����^� 3�^� ������Vh(�h�   hD �����������t���   ��t�t$����^� 3�^� ������Vh(�h�   hD ����������t���   ��t�t$����^� 3�^� ������Vh(�h�   hD ���I�������t���   ��t��^��3�^����������������Vh(�h�   hD ���	�������t���   ��t�t$���t$�t$��^� 3�^� ��������������Vh(�h�   hD ����������t���   ��t�t$����^� ������������Vh(�h�   hD ���y�������t���   ��t�t$���t$�t$��^� 3�^� ��������������Vh(�h�   hD ���)�������t���   ��t��^��3�^����������������h(�jhD ���������t	�@��t��3��������������j�h�yd�    P��VW�P�3�P�D$ d�    h(�h�   hD �D$    ��������u)� ��t$0�HV�I�у��ƋL$ d�    Y_^�� ��t$4���   �L$Q�Ћ�� ��|$8�IW�I�D$4   �ѡ �W�@V�@�Ћ ��D$$�IP�I�D$$   �D$@ �у��ǋL$ d�    Y_^�� ������������h(��t$hD ����������������̡ ����   �AP���   ��Y�������̡ ��t$�@8Q�@D�Ѓ�� �������̡ ��@8�@<����̡ �V�@8�t$�@@�6�Ѓ��    ^���t$� ��t$�@8�t$�@�t$�t$�t$Q�Ѓ�� �����t$� ��t$�@8�t$�@�t$�t$Q�Ѓ�� �������̡ ��@8� �����̡ �V�@8�t$�@�6�Ѓ��    ^���t$� ��t$�@8�t$�@Q�Ѓ�� � ��t$�@8�t$�@Q�Ѓ�� ���̡ �Q�@8�@�Ѓ���������������̡ ��t$�@8Q�@ �Ѓ�� ���������t$� ��t$�@8�t$�@$�t$�t$Q�Ѓ�� �������̡ ��t$�@8�t$�@(Q�Ѓ�� �����t$� ��t$�@8�t$�@,Q�Ѓ�� �t$� ��t$�@8�t$�@Q�Ѓ�� � ��t$�@8�t$�@0Q�Ѓ�� �����t$� ��t$�@8�t$�@4Q�Ѓ�� � ��t$�@8Q�@8�Ѓ�� �������̋L$� ��P�APP�A@P�A0P�A P�AP���   Q�t$�Ѓ����������������̡ ��@���   �� ��@���  �� ��@�@,����̡ ��@���  ��j�h�yd�    PQV�P�3�P�D$d�    �D$    � ��t$�@V�@�D$    �Ћ �V�I�D$    �I8�D$   �у��ƋL$d�    Y^���������̡ ��@�@<����̡ ��@�@@����̡ ��@�@D����̡ ��@�@H����̡ ��@�@L����̡ ��@�@P����̡ ��@��<  �� ��@��,  ���t$� ��t$�@�t$���   �t$�t$h�6  �Ѓ����̡ ��@�@�����j�h zd�    P�� �P�3�P�D$$d�    � ��L$�@Q�@�С �j �@j��@�L$hd�Q���t$H�D$P�D$0P�D$L    ������ ��L$$�@Q�@�D$P�С ��L$8�@Q�@�С ��L$<�@Q�@�D$X�����Ѓ�,�L$$d�    Y��,���������������̡ ��@���  �� ��@��8  ��j�h\zd�    P��VW�P�3�P�D$ d�    �D$    � ��L$�@Q��  �Ћ�� ��|$4�IW�I�D$0   �ѡ �W�@V�@�Ћ ��D$ �IP�I�D$    �D$< �у��ǋL$ d�    Y_^�� ������������j�h�zd�    P��VW�P�3�P�D$ d�    �D$    � ��L$�@Q��  �Ћ�� ��|$4�IW�I�D$0   �ѡ �W�@V�@�Ћ ��D$ �IP�I�D$    �D$< �у��ǋL$ d�    Y_^�� �����������̡ ��@��x  �� ��@��|  �� ��@���  �� ��@���  �� ��@���  �� ��@�@T����̡ ��@�@X����̡ ��@�@\����̡ ��@�@`����̡ ��@���  �� ��@�@d����̡ ��@�@h����̡ ��@�@l����̡ ��@�@p����̡ ��@�@t����̡ ��@��D  �� ��@��  �� ��@�@x����̡ ��@��@  ��j�h�zd�    PQV�P�3�P�D$d�    �D$    �t$���D$    �3���� �V�I�t$$�I|�D$    �D$   �у��ƋL$d�    Y^������������̡ ��@���   �� ��@��d  �� ��@��h  �� ��@���  �� ��@���   ��j�h�zd�    PQV�P�3�P�D$d�    �D$    �t$���D$    ��'��� �V�I�D$    ���   �D$   �у��ƋL$d�    Y^�������������̡ ��@��`  �� ��@��  �� ����@�t$ ���   �L$Q�ЋL$$�~ f��~@f�A�~@f�A���� ��������������̡ ��@���  ���t$�D$� ����@�D$�D$���   �$�t$�Ѓ�����������̡ ��@���   �� ��@���   �� ��@���  �� ��@���  �� ��@��   �� ��@��  �� ��@��l  �� ��@���  �� ��@���  �� ��@���  �� ��@���  �� ��@���  �� ��@���  ��j�h4{d�    P��VW�P�3�P�D$ d�    �t$4�D$    � ��L$�@Q���  �Ћ�� ��|$8�IW�I�D$4   �ѡ �W�@V�@�Ћ ��D$$�IP�I�D$$   �D$@ �у��ǋL$ d�    Y_^�� ��������j�hp{d�    P��VW�P�3�P�D$ d�    �t$4�D$    � ��L$�@Q���  �Ћ�� ��|$8�IW�I�D$4   �ѡ �W�@V�@�Ћ ��D$$�IP�I�D$$   �D$@ �у��ǋL$ d�    Y_^�� �������̡ ��@���  �� ��@���  ����� ��T$�@R���   �T$R�T$RQ�����#D$���̃�� ��T$�@R���   �T$R�T$RQ�����#D$���̃�� ��$�@R���   �T$R�T$RQ�����#D$����̡ ��@���   �� ��@���   �� ��@���   �� ��@���   �� ��@���   �� ��@���   �� ��@��  �� ��@��\  ��j�h�{d�    P�� �P�3�P�D$$d�    �t$8�D$    � ��L$�@Q��t  �Ѓ��t$4���D$0   �V����L$�D$   �D$, 耹���D$4�L$$d�    Y��,������������̡ ��@��H  �� ��@��T  �� ��@��p  �� ��@��8  ����  �P�3ĉ�$   ��$  P��$  �D$h   P�L�����x	=�  |'�� �hh��@hH  ��0  �Ѓ�Ƅ$�   � ��$�@Q��4  h`��Ћ�$  ��3��NG  ��  �������������������������t$$�D$�t$$�P�t$$� ��t$$�@0�t$$���   �t$$�t$$�t$$RQ�Ѓ�(�$ ��t$$�D$�t$$�P�t$$� ��t$$�@0�t$$���   �t$$�t$$�t$$RQ�Ѓ�(�$ ��t$$� ��t$$�@0�t$$���   �t$$�t$$�t$$�t$$�t$$�t$$Q�Ѓ�(�$ ����̡ �Q�@0���   �Ѓ������������̡ ��t$�@0�t$���   Q�Ѓ�� ��t$� ��t$�@0�t$���   �t$Q�Ѓ�� ��������̡ �Q�@0���   �Ѓ��������������t$� ��t$�@0�t$���   �t$Q�Ѓ�� ��������̡ ��@0���   �� �V�@0�t$���   �6�Ѓ��    ^���������������j�h�{d�    P��V�P�3�P�D$d�    �t$8�D$    � ��t$8�@�t$8��X  �L$Q�ЋЋt$<j �    �F    � �R���   V�@�D$@   �Ћ ��D$(���   P�	�D$(   �D$D �у� �ƋL$d�    Y^�� ������������j�h(|d�    P��(V�P�3�P�D$0d�    hLGOg�L$ �D$    �F��j P�D$hicMCP�D$H   ��������L$�D$8�[��� ��L$���   Q�@T�Ѓ���u�L$@�����"� ��L$���   Q�@T�ЋL$D��P����� ��D$���   P�	�D$   �D$< �ыD$D���L$0d�    Y^��4��������̡ ��@���  �� ��@���  �� ��@���  ��j�hd|d�    P��VW�P�3�P�D$ d�    j �t$D�D$    �t$D� ��t$D�@�t$D��t  �L$$Q�Ћ�� ��|$H�IW�I�D$D   �ѡ �W�@V�@�Ћ ��D$4�IP�I�D$4   �D$P �у�(�ǋL$ d�    Y_^�� ����������j�h�|d�    P��V�P�3�P�D$d�    �t$<�D$    �t$<� ��t$<�@�t$<���  �L$Q�ЋЋt$@j �    �F    � �R���   V�@�D$D   �Ћ ��D$,���   P�	�D$,   �D$H �у�$�ƋL$d�    Y^�� ��������j�h�|d�    P��$�P�3�P�D$(d�    � ��@��p  �Ѕ���   h���L$���� ��t$8�@h���@4�L$�D$8    �С ��t$<�@h���@4�L$��j �D$P�D$hicMCP����� ��L$���   Q� �Ѓ��L$�D$0�����]���L$(d�    Y��0��������������j�h}d�    P��(VW�P�3�P�D$4d�    �D$    � ��@��p  �Ѕ�u)� ��t$D�HV�I�у��ƋL$4d�    Y_^��4�h!���L$$���� ��t$H�@h!���@4�L$(�D$D   ��j �D$$P�D$hicMCP����P� ��D$P���   �@H�Ћ ��|$X�IW�I���ы �W�AV�@�Ћ ��D$0���   P�	�D$0   �D$`�у�$�L$ �D$< �!���ǋL$4d�    Y_^��4��������������j�hK}d�    P��(VW�P�3�P�D$4d�    �D$    � ��@��p  �Ѕ�u)� ��t$D�HV�I�у��ƋL$4d�    Y_^��4�h����L$$�H��� ��t$H�@h����@4�L$(�D$D   ��j �D$$P�D$hicMCP�����P� ��D$P���   �@H�Ћ ��|$X�IW�I���ы �W�AV�@�Ћ ��D$0���   P�	�D$0   �D$`�у�$�L$ �D$< �����ǋL$4d�    Y_^��4��������������j�hv}d�    P��$V�P�3�P�D$,d�    � ��@��p  �Ѕ�u�L$,d�    Y^��0�h#���L$�)��� ��t$<�@h#���@4�L$ �D$<    ��j �D$P�D$hicMCP����P� ��D$H���   �@8�Ћ ������   �D$�	P�D$L �у��L$�D$4���������ƋL$,d�    Y^��0��������j�h�}d�    P��$V�P�3�P�D$,d�    � ��@��p  �Ѕ�u�L$,d�    Y^��0�hs���L$�9��� ��t$<�@hs���@4�L$ �D$<    ��j �D$P�D$hicMCP�����P� ��D$H���   �@8�Ћ ������   �D$�	P�D$L �у��L$�D$4���������ƋL$,d�    Y^��0�������̡ ��@���  �� ��@���  �� ��@��@  ��V�t$���t� �Q�@��D  �Ѓ��    ^���������̡ ��@��H  �� ��@��L  �� ��@��P  �� ��@��T  �� ��@��X  �� ��@��\  �� ��@��d  �� ��@��h  �� ��@��l  �� ��@���  �� ��@���  �� ��@���  �� ��@��P  �� ��@���  ��j�h�}d�    P���P�3�P�D$d�    �t$0�D$    � ��L$�@Q���  �Ѓ��L$,P�D$(   �'���L$�D$   �D$$ �1���D$,�L$d�    Y��$�������������̡ ��@���  �� ��@���  �� ��@���  �� ��@���  �� ��@���  �� ��@���  �� ��@��l  �� ��@���  �� ��@���  �� ��@��$  �� ��@��(  �� ��@��,  �� ��@��0  �� ��@��<  �� ��@��  �� ��@��`  �� ��@��\  ��h8�jh�f �Ϥ������t	�@��t�����������������j�h~d�    PQV�P�3�P�D$d�    h8�jh�f �D$     �u���������t9�~ t3�t$L�D$$�t$L�t$L�t$L�t$L����P�����t$L�F�Ѓ�4�������L$ �D$�����o����ƋL$d�    Y^���������������h8�jh�f ��������t	�@��t��3��������������h8�jh�f 迣������t	�@��t��3��������������h8��t$h�f 荣�������������̃� �(�V���.�vf(�fT`�f/�f(�fT`��T$�L$�L$�-  f/��#  �8�f/�vFf/�v@�,��,���   ��$    ������ʅ�u�fn�����^��^��.�v^�� �f/�v(��(��H��^��%��f/�v4(��Y��Y��Y��D$(��Y��.�v(��L$�L$f/�v(��D$�D$�f��D$�D$�i<  �\$�D$f/0��L$�L$�D$�D$s���^���F�^��F^�� �W������F^�� �����������������D$�@�f/�V��w�P�f/�v(��Yؖ���X0��D$�D$�$�;  �ؖ������F�������^� ���̃��L$�T$3�W�f/�fT`��X0���3�f/�V����3��L$�D$;������$�L$�);  ��D$ fT`��D$ �X0��D$ �D$ �$��:  ����\$ �D$ ��f/��Fv'� �h���@j��0  ��������F�|$ u�fWp����������^��� ������������D$���f/�V���Fv'� �hԗ�@j,��0  ��������F^� ���������U�����M�����<f/�V��v'� �h���@j5��0  ��������M��Y����D$8�D$8�$��9  �\$8�F�$�9  �D$8�\$@�^D$@�D$@�D$@�$�9  ��E�$�9  ���^�������^��]� ����������̋L$��`������̋L$��`�������V��h�*����F    � �V�@Ph�'� h�'�Ѓ��F��^����������̃y ���u� ��q�@P�@��Y��̋I��u3�� � �j �t$�@P�t$�@Q�Ѓ�� �����̋I��t� ��t$�@PQ�@�Ѓ�� ̋I��t� ��t$�@PQ�@�Ѓ�� ��    �A    ���V����t&� �Q�@P�@L�С ��6�@P�@<�Ѓ��    ^����������������SUVW�����t� �Q�@P�@<�Ѓ��    �G    �\$�l$h�*S�o� �h�'�@Ph�'�@8U�t$(�Ѓ�3����~D���x u�@   � ��HP���p�A�Ѓ�� �V�@P�7�@@�Ћ�F���A;�|�3�9_^]��[� �������������t$�D$�t$�p�,���� ���������SVW��3�9w~>�\$� �V�@P�7�@@�ЋЃ���t,� �j �APS�@jR�Ѓ���tF;w|�_^�   [� � ��7�@P�@L�Ѓ�3�_^[� ̡ ��1�@P�@D�Ѓ��������������̡ ��1�@P�@H��Y���������������̡ ��1�@P�@L��Y���������������̡ ��@P�@P����̡ ��@P�@T����̡ ��@P���   �� ��@P���   ���L$��`�������V��~ ���u� ��v�@P�@�Ѓ��D$t	V�!�������^� ��������3��������������̡ �Q�@L���   �Ѓ������������̡ ��t$�@L�t$���   Q�Ѓ�� ̡ �V�@L�񋀠   V�Ћȡ �����u�@LQ�t$���   V�Ѓ�^� ���   �@P�Ћ �P���   �L$�BH��^� ̡ �Q�@L��(  �Ѓ������������̡ ��t$�@L�t$��,  Q�Ѓ�� ̡ ��@L� �����̡ �V�@@�t$�@�6�Ѓ��    ^�̡ ��@L���   �� �V�@@�t$�@�6�Ѓ��    ^��j�hM~d�    P���P�3�P�D$d�    �t$0�D$    � �Q�@L�L$�@Q�Ѓ��L$,P�D$(   �9
���L$�D$   �D$$ �C
���D$,�L$d�    Y��$� ������������̡ ��t$�@L�t$�@Q�Ѓ�� ���̡ ��t$�@LQ���   �Ѓ�� ����̡ �Q�@L�@�Ѓ���������������̡ �Q�@L�@�Ѓ���������������̡ �Q�@L�@�Ѓ�����������������t$� ��t$�@L�t$�@ Q�Ѓ�� � ��t$�@LQ��4  �Ѓ�� ������t$� ��t$�@L�t$�@$Q�Ѓ�� �t$� ��t$�@L�t$�@(�t$Q�Ѓ�� �����������̡ �Q�@L�@,�Ѓ���������������̡ �Q�@L�@0�Ѓ���������������̡ �Q�@L�@4�Ѓ���������������̡ �j �@LQ�@8�Ѓ�������������̡ ��t$�@L�t$��  Q�Ѓ�� ̡ ��@L���   �� ��@L���   �� ��@L��l  �� ��@L���   �� ��@L���   �� ��@L���   �� ��@L���   �� ��@L���   �� ��@L���   �� ��t$�@LQ�@<�Ѓ�� �������̡ ��@L���   �� �Q�@L�@��Yá ��t$�@L�t$�@@Q�Ѓ�� ���̡ �j �@L�t$�@DQ�Ѓ�� �����̡ �j�@L�t$�@DQ�Ѓ�� �����̡ �j �@L�t$�@HQ�Ѓ�� �����̡ �j�@L�t$�@HQ�Ѓ�� �����̡ �Q�@L���   �Ѓ�������������j�h�~d�    P���P�3�P�D$d�    �t$0�D$    � �Q�@L�L$��  Q�Ѓ��L$,P�D$(   �F���L$�D$   �D$$ �P���D$,�L$d�    Y��$� ����������j�h�~d�    P��$SV�P�3�P�D$0d�    ���D$     �D$(    �D$P�L$�D$<    �D$�  �D$    �D$     ����j �D$$P�D$P���D$D�$  ���L$���D$8 ������t3��� ��L$ ���   Q�@8�Ѓ���� ��D$ ���   P�	�D$<�����у��ƋL$0d�    Y^[��0�����������j�h�~d�    P��$V�P�3�P�D$,d�    ���D$   �D$$   �D$P�L$�D$8    �D$�  �D$    �D$    �,���j�D$ P�D$P���D$@��#  �L$�D$4 ����� ��L$���   Q� �D$8�����Ѓ��L$,d�    Y^��0�������j�hd�    P��(SV�P�3�P�D$4d�    ���D$    �D$$    �D$,    �D$P�L$�D$@   �D$�  �D$     �D$$    �c���j �D$(P�D$P���D$H��"  ���L$���D$<�������t�L$D�����"� ��L$$���   Q�@L�ЋL$H��P�g���� ��D$$���   P�	�D$   �D$@ �ыD$H���L$4d�    Y^[��4� ����������j�hcd�    P��(SV�P�3�P�D$4d�    ���D$    �D$$    �D$,    �D$P�L$�D$@   �D$�  �D$     �D$$    �S���j �D$(P�D$P���D$H��!  ���L$���D$<������t�L$D�����"� ��L$$���   Q�@L�ЋL$H��P�W���� ��D$$���   P�	�D$   �D$@ �ыD$H���L$4d�    Y^[��4� ����������j�h�d�    P��$V�P�3�P�D$,d�    �� ��t$<�D$     �D$(    ���   �L$ �@(Q�Ѓ��D$P�L$�D$8    �D$�  �D$    �D$    �0���j�D$ P�D$P���D$@��   �L$�D$4 蚿��� ��L$���   Q� �D$8�����Ѓ��L$,d�    Y^��0� ��������j�h�d�    P��$V�P�3�P�D$,d�    �� ��t$<�D$     �D$(    ���   �L$ �@(Q�Ѓ��D$P�L$�D$8    �D$�  �D$    �D$    �P���j�D$ P�D$P���D$@��  �L$�D$4 躾��� ��L$���   Q� �D$8�����Ѓ��L$,d�    Y^��0� ��������j�h�d�    P��,SV�P�3�P�D$8d�    ���D$(    �D$0    �D$P�L$�D$D    �D$ �  �D$$    �D$(    苼��j �D$,P�D$P���D$L�#  ���L$���D$@ ������tW��D$�D$�� ��L$(���   Q�@<�Ѓ�� ��\$�L$(���   Q� �D$D�������D$���L$8d�    Y^[��8�������������j�h�d�    P��V�P�3�P�D$$d�    ���D$4�D$   �D$�D$P�L$8�D$0    �D$�  �D$    �D$    舻��j�D$P�D$<P���D$8�0  �L$4�D$, ����� ��L$���   Q� �D$0�����Ѓ��L$$d�    Y^��(� j�h:�d�    P��$SV�P�3�P�D$0d�    ���D$     �D$(    �D$P�L$�D$<    �D$�  �D$    �D$     �˺��j �D$$P�D$P���D$D�c  ���L$���D$8 �0�����t3��� ��L$ ���   Q�@8�Ѓ���� ��D$ ���   P�	�D$<�����у��ƋL$0d�    Y^[��0�����������j�he�d�    P��$V�P�3�P�D$,d�    ��D$<�D$   �D$$�D$P�L$�D$8    �D$�  �D$    �D$    �ܹ��j�D$ P�D$P���D$@�  �L$�D$4 �F���� ��L$���   Q� �D$8�����Ѓ��L$,d�    Y^��0� ����j�h��d�    P��$SV�P�3�P�D$0d�    ���D$     �D$(    �D$P�L$�D$<    �D$�  �D$    �D$     ����j �D$$P�D$P���D$D�  ���L$���D$8 耺����t:� ��t$@���   W��	�����D$ P�F�D$<�����у��K� ��L$ ���   Q�@P���~ �t$D� �f��~@���   �D$$�	Pf�F�D$@�����у��ƋL$0d�    Y^[��0� �j�h��d�    P��$V�P�3�P�D$,d�    �� ��t$<�D$     �D$(    ���   �L$ �@,Q�Ѓ��D$P�L$�D$8    �D$�  �D$    �D$    �з��j�D$ P�D$P���D$@�x  �L$�D$4 �:���� ��L$���   Q� �D$8�����Ѓ��L$,d�    Y^��0� ��������j�h�d�    P��$SV�P�3�P�D$0d�    ���D$     �D$(    �D$P�L$�D$<    �D$�  �D$    �D$     ����j �D$$P�D$P���D$D�  ���L$���D$8 �p�����t:� ��t$@���   W��	�����D$ P�F�D$<�����у��K� ��L$ ���   Q�@P���~ �t$D� �f��~@���   �D$$�	Pf�F�D$@�����у��ƋL$0d�    Y^[��0� �j�h�d�    P��$V�P�3�P�D$,d�    �� ��t$<�D$     �D$(    ���   �L$ �@,Q�Ѓ��D$P�L$�D$8    �D$�  �D$    �D$    �����j�D$ P�D$P���D$@�h  �L$�D$4 �*���� ��L$���   Q� �D$8�����Ѓ��L$,d�    Y^��0� �������̡ ����@Lj�t$���   Q�L$Q�ЋL$$�~ f��~@f�A���� � ��̡ ����@Lj �t$���   Q�L$Q�ЋL$$�~ f��~@f�A���� � ���j�h<�d�    P��$SV�P�3�P�D$0d�    ���D$     �D$(    �D$P�L$�D$<    �D$�  �D$    �D$     �{���j �D$$P�D$P���D$D�  ���L$���D$8 ������t:� ��t$@���   W��	�����D$ P�F�D$<�����у��K� ��L$ ���   Q�@P���~ �t$D� �f��~@���   �D$$�	Pf�F�D$@�����у��ƋL$0d�    Y^[��0� �j�hg�d�    P��$V�P�3�P�D$,d�    �� ��t$<�D$     �D$(    ���   �L$ �@,Q�Ѓ��D$P�L$�D$8    �D$�  �D$    �D$    �0���j�D$ P�D$P���D$@��  �L$�D$4 蚴��� ��L$���   Q� �D$8�����Ѓ��L$,d�    Y^��0� ��������j�h��d�    P��$SV�P�3�P�D$0d�    ���D$     �D$(    �D$P�L$�D$<    �D$�  �D$    �D$     �k���j �D$$P�D$P���D$D�  ���L$���D$8 �г����t:� ��t$@���   W��	�����D$ P�F�D$<�����у��K� ��L$ ���   Q�@P���~ �t$D� �f��~@���   �D$$�	Pf�F�D$@�����у��ƋL$0d�    Y^[��0� �j�h��d�    P��$V�P�3�P�D$,d�    �� ��t$<�D$     �D$(    ���   �L$ �@,Q�Ѓ��D$P�L$�D$8    �D$�  �D$    �D$    � ���j�D$ P�D$P���D$@��  �L$�D$4 芲��� ��L$���   Q� �D$8�����Ѓ��L$,d�    Y^��0� ��������j�h�d�    P��$SV�P�3�P�D$0d�    ���D$     �D$(    �D$P�L$�D$<    �D$�  �D$    �D$     �[���j �D$$P�D$P���D$D��  ���L$���D$8 �������t3��� ��L$ ���   Q�@8�Ѓ���� ��D$ ���   P�	�D$<�����у��ƋL$0d�    Y^[��0�����������j�h�d�    P��$V�P�3�P�D$,d�    ��D$<�D$   �D$$�D$P�L$�D$8    �D$�  �D$    �D$    �l���j�D$ P�D$P���D$@�  �L$�D$4 �ְ��� ��L$���   Q� �D$8�����Ѓ��L$,d�    Y^��0� ����j�h>�d�    P��$SV�P�3�P�D$0d�    ���D$     �D$(    �D$P�L$�D$<    �D$�  �D$    �D$     諮��j �D$$P�D$P���D$D�C  ���L$���D$8 ������t:� ��t$@���   W��	�����D$ P�F�D$<�����у��K� ��L$ ���   Q�@P���~ �t$D� �f��~@���   �D$$�	Pf�F�D$@�����у��ƋL$0d�    Y^[��0� �j�hi�d�    P��$V�P�3�P�D$,d�    �� ��t$<�D$     �D$(    ���   �L$ �@,Q�Ѓ��D$P�L$�D$8    �D$�  �D$    �D$    �`���j�D$ P�D$P���D$@�  �L$�D$4 �ʮ��� ��L$���   Q� �D$8�����Ѓ��L$,d�    Y^��0� ��������j�h��d�    P��$SV�P�3�P�D$0d�    ���D$     �D$(    �D$P�L$�D$<    �D$�  �D$    �D$     蛬��j �D$$P�D$P���D$D�3  ���L$���D$8 � �����t3��� ��L$ ���   Q�@8�Ѓ���� ��D$ ���   P�	�D$<�����у��ƋL$0d�    Y^[��0�����������j�h��d�    P��$V�P�3�P�D$,d�    ��D$<�D$   �D$$�D$P�L$�D$8    �D$�  �D$    �D$    謫��j�D$ P�D$P���D$@�T  �L$�D$4 ����� ��L$���   Q� �D$8�����Ѓ��L$,d�    Y^��0� ����j�h�d�    P��$SV�P�3�P�D$0d�    ���D$     �D$(    �D$P�L$�D$<    �D$�  �D$    �D$     ����j �D$$P�D$P���D$D�  ���L$���D$8 �P�����t3��� ��L$ ���   Q�@8�Ѓ���� ��D$ ���   P�	�D$<�����у��ƋL$0d�    Y^[��0�����������j�h�d�    P��$V�P�3�P�D$,d�    ��D$<�D$   �D$$�D$P�L$�D$8    �D$�  �D$    �D$    �����h�   �D$ P�D$P���D$@�  �L$�D$4 �c���� ��L$���   Q� �D$8�����Ѓ��L$,d�    Y^��0� �������t��t��t3�ø   ���̡ �Q�@L�@L�Ѓ���������������̡ �Q�@L�@P�Ѓ�����������������t$� ��t$�@L�t$���  Q�Ѓ�� ������������̡ ��t$�@LQ��  �Ѓ�� ����̡ ��t$�@LQ���   �Ѓ�� ����̡ �Q�@L�@X�Ѓ�����������������t$� ��t$�@L�t$�@\Q�Ѓ�� j�h@�d�    P��0SVW�P�3�P�D$@d�    �� ��@L�@�Ћ؅�u�L$@d�    Y_^[��<� �L$�����D$H    �D$(    �D$0    �D$4    �D$<    �D$8    �t$P�D$�D$0� ��\$(�@h]  �@0�L$�D$P�С �j ���   j �@S���Ѕ���   � �S�@L�@�Ћ�������   ��� ����   �΋R(�ҋ��D$$Ph�   �t$0���������ts�L$<��tk� �j ���   ���   �ЋЅ�tP� �V���   �ʋ@<�С ��L$<���   Q���   �Ѓ���t� �V�@@�@�Ѓ������`����+� �S�@@�@�С ��L$@���   Q���   �Ѓ�3ۍL$$�D$H 蕹���L$�D$H�����d����ËL$@d�    Y_^[��<� ������������̡ �Q�@L�@`�Ѓ���������������̡ �Q�@L�@d�Ѓ���������������̡ ��t$�@LQ�@h�Ѓ�� �������̡ �Q�@L��D  �Ѓ������������̡ �Q�@L�@l�Ѓ���������������̡ ��t$�@LQ���   �Ѓ�� ����̡ ��@L�@����̡ �V�@@�t$�@�6�Ѓ��    ^�̡ �Q�@L���   ��Y�������������̡ �Q�@L���   �Ѓ��������������t$� ��t$�@L�t$���   �t$�t$Q�Ѓ�� ������t$� ��t$�@L�t$���   Q�Ѓ�� ��������������t$� ��t$�@L�t$��   �t$Q�Ѓ�� ����������t$� ��t$�@L�t$��   Q�Ѓ�� ������������̡ ��@L��H  �� ��@L��L  �� ��@L��P  �� ��@L��T  �� ��@L��p  �� ��@L��t  �� ��@L���  �� ��@L���  �� ��@L���  �� ��@L���  ���T$ V�t$�D$h�Sh�Sh�Sh�SR�t$4�q�t$4�Q�t$4� ����@L�$�t$4���   VQ�Ѓ�4^�  ����̡ ��@���   �� ��@���   �� ��@���   �� ��@���   �� ��@���   �� �V�@�t$���   �6�Ѓ��    ^��������������̡ �V�@L�@�Ћ���u^á �j �t$�@�t$��h  �t$V�Ѓ���u� �V�@@�@�Ѓ�3���^�������������̡ �j �H�t$�D$�� P�t$��h  �t$�Ѓ�������̡ ��@���   �� ��@L���   ���t$� ��t$�@�t$���   �t$ �t$ �t$ �t$�Ѓ��j�hk�d�    P�� V�P�3�P�D$(d�    �D$    �D$    �D$    �D$    �D$    �D$$    �D$     � ��D$0    ���   ���   �ЉD$�t$8�D$0��t<��t8� �j�QLP���   ���ЋD$�D$ �D$Ph=���t$����������   � ��L$���   Q���   �D$4 �Ѓ��L$�D$    �D$0���������ƋL$(d�    Y^��,������������j�h��d�    P�� V�P�3�P�D$(d�    �D$    �D$    �D$    �D$    �D$    �D$$    �D$     � ��D$0    ���   ���   �ЉD$�t$8�D$0��t<��t8� �j�QLP���   ���ЋD$�D$ �D$Ph<���t$�Ӻ��������   � ��L$���   Q���   �D$4 �Ѓ��L$�D$    �D$0���������ƋL$(d�    Y^��,�����������̡ ��@L���   �� ��@L���   �� ��@L��  �� ��@L��@  ���L$�� �������̋L$�t$��P��̋L$�t$��t$�P����������������t$�L$�t$��t$�t$�P������̡ �V���   �񋀌   V�Ѓ��    ^��������������̋D$HV����   �$�U�   ^áL�@�L���uU�t$�v����=�6  }�����^Ët$��t�jh��jmj���������t	���v���3��H���tV���~}���   ^��t$�t$�Z����������H^�^�'����L�u.�*����%����5H���t���Dx��V�������H�    �   ^Ã��^ÐMT�T�TFTU�T�������������L$u�D$�@��D$�D��   � �A    �    �A    �A   ������t$� ��t$�@@�t$�@Q�Ѓ�� � ��t$�@@Q�@�Ѓ�� �������̡ ��t$�@@�t$�@Q�Ѓ�� ���̡ ��t$�@@Q�@ �Ѓ�� �������̡ ����   �@�� ����   �@�� ����   �@ �� ����   �@$�� ����   ���   ��������������̡ ����   ��D  ��������������̡ ��t$�@@Q�@L�Ѓ�� �������̡ �Q�@@�@H�Ѓ���������������̡ ����   ���   ��������������̡ ����   ���   ��������������̡ �Q�@H���   �Ѓ�������������V��L$��t2�T$� ����   ��t
�@@R��^� �T$�@D��tR��^� V��^� ��������������̡ ��@@�@0�����V�t$���t� �Q�@@�@�Ѓ��    ^������������̡ �V�@@��@V�ЋЋD$����t��#��С �R�@@V�@�Ѓ�^� �����t$�D$� ������   �$�t$���   �t$�t$�t$��� �������̡ ����   ���   ��������������̡ �Q�@H���   �Ѓ������������̡ ��t$�@HQ��d  �Ѓ�� ����̡ ��@@�@T����̡ ��@@�@X����̡ ��@@�@\����̡ ��@@�@`����̡ ��@@�@d����̡ ��@@�@h����̡ ��@@�@l����̡ ��@@���   �� ��@@�@t����̡ ��@@�@x����̡ ��@@�@|����̡ ��@@���   �� ��@@���   �� ��@@���   �� ����   �@t�� ��@@���   �� ��@@���   �� ��@@���   �� ��@@���   �� ��@@���   �� ��@@���   �� ��@@���   ��V�t$���t� �Q�@@�@�Ѓ��    ^������������̡ ��@@�@0����̡ �j�@@�L$�@4Qj �Ѓ�������̡ �j�@@�L$�@4Qh   @�Ѓ����̡ ��t$�@@�t$�@4j �Ѓ������̡ ��@|� ������V�t$���t� �Q�@|�@�Ѓ��    ^������������̡ ��@|�@ �����V�t$���t� �Q�@|�@(�Ѓ��    ^������������̡ ��@ �@H����́|$qF uKW�|$��tA� ��t$���   �ϋ@D�С ��t$�@@�@,�Ћ ����ЋAW�t$�@p����_����������̡ ��@��T  �� �S�@@V�@,W�t$�Ћ ��t$�I@�؋I,�ы ����yh��hE  �ˋ��)���Ph��hE  ������P��T  �Ѓ�_^[���%��;P�u���:  ��%|��%x�U���EV��t%Whc�~��7jV�  �EtW�����Y��_��  �EtV����Y��^]� Vh�   �,�Y��V����������u3�@^Ã& �t  h+e�>  �$Xe�2  Y3�^�U��QQ�} SVW�)  �T����  H�T�d�   3��P�}�����;�t3�������u���E�   �=��tj�  Y�  �5�������u����   �5�����؉u�]��;�r\9;t�W��9t��3��W��������5���5����5���E��֋M�9Mu�u9Et���M�u�E��띃��tV�t�YW������������=��9}���   3���   3��   �}��   d�   3��P������;�t3�������u��3�F9=��j_t	j��  �5h��h�����   �  YY��u�h��h����  Y�=��Y��u3���=�� th����  Y��t�uW�u����T�3�@_^[�� U��}u�  �u�u�u�   ��]� jh���  3�@���u�3ۉ]��}�=`��E���u9=T���   ;�t��u8����t�uW�u�Ћ��u����   �uW�u�������u����   �uW�u��������u��u.��u*�uS�u������uS�u�@�������t	�uS�u�Ѕ�t��uK�uW�u�������#��u�t4����t+�uW�u�Ћ���M�� �E�QP�K  YYËe�3ۋ�u�]��E������   ����  Ëu��`������̃=�� t3��Vjj �@�YY��V����������ujX^Ã& 3�^�jh ��*  �5���5��։E���u�u�H�Y�ej�}  Y�e� �5���։E��5���։E��E�P�E�P�u�5���P�U  �����}��u��֣���u��֣���E������   ����  Ë}�j�  Y�U���u�P��������YH]��������������%l��%h�U����j�t���  �u��  �=t� YYuj��  Yh	 ���  Y]�U���$  j��  ��tjY�)�X��T��P��L��5H��=D�f�p�f�d�f�@�f�<�f�%8�f�-4���h��E �\��E�`��E�l����������  �`��d��X�	 ��\�   �h�   jXk� ǀl�   jXk� �P��L�jX�� �T��L�h��������jh@��"  �e� �]�Ë}�ǋu��u�e� O�}x+�u���U��3�@�E��E������   �#  � �}�]�u�E��u�uWSV�   �jh`��  �e� �Mx:�M+M�M�U��E�E�E� �E��E��8csm�t�E�    �E���  �e��E������  � ��%D��%$��%(���������������U��ES�H<�V�A�Y��3��W��t�}�p;�r	�H�;�r
B��(;�r�3�_^[]��������������U��j�h��h�ed�    P��SVW�P�1E�3�P�E�d�    �e��E�    h   �|   ����tT�E-   Ph   �R�������t:�@$���Ѓ��E������M�d�    Y_^[��]ËE� 3Ɂ8  �����Ëe��E�����3��M�d�    Y_^[��]�������U��E�MZ  f9t3�]ËH<�3��9PE  u�  f9Q��]�U����P��e� �e� VW�N�@��  ��;�t��t	�УT��f�E�P���E�3E�E�� �1E���1E��E�P���M�3M�E�3M�3�;�u�O�@����u��G  ��ȉP��щT�_^��VW�$��$�����t�Ѓ�;�r�_^�VW�,��,�����t�Ѓ�;�r�_^���%0��%4�hx��   Y�������������h�ed�5    �D$�l$�l$+�SVW�P�1E�3�P�e��u��E��E������E��E�d�    ËM�d�    Y__^[��]Q�U���u�u�u�uh \hP��5   ��]��%8��%<��%���%P��%T��%X��%\��%`��%d��%��������̍M������M�� ����T$�B�J�3�������������M������M������T$�BԋJ�3������ԟ�����M�������T$�B��J�3��a�������g����M��ϰ���M������M�鿰���M������M�鯰���M������M�韰���M��w���h<�h5  hP��E�P蟰����ÍM��s����T$�B؋J�3���������������������̋M����%����M������T$�B�J�3������@������̋M��(����T$�B��J�3������ܠ�����������������h0�h  hP��E�P�������ËM��ܯ���T$�B�J�3��;������A���̋E����   �e���M�X���ÍM��o����M���d����T$�B�J�3����������������������̍M�������T$�B؋J�3�������t������������������̍M���d���T$�B��J�3������������hx�j;hP��E�P������ËT$�B��J�3��c�������i����M��Ѯ���M��ɮ���EЃ��   �e���M鱮��ËT$�BЋJ�3������`��%����M�鍮���M�酮���EЃ��   �e���M�m���ÍM��d����T$�BЋJ�3�������<�������M��A����M��9����EЃ��   �e���M�!���ÍM������M������T$�BЋJ�3������������M������M������EЃ��   �e���M�ͭ��ÍM��ĭ���M�鼭���M�鴭���T$�BЋJ�3��#�������)����M�鑭���E����   �e���M��y���ËE����   �e���M��`���ËT$�B��J�3�������С������M��<����E����   �e���M��$���ËE����   �e���M�����ËT$�B��J�3��y������������������������̍M��ج���E����   �e���M�����ËT$�B�J�3��.����4��4������̍M��Xb���Eԃ�t�e���M�Db��ËT$�B��J�3�������h�������������̍�h����b����X����J����M��b���M���a���M���a���M���a���T$��\�����X���3��������������������̍M�������E����   �e���M����ËT$�B�J�3��N������T����M�霫���T$�B�J�3��+������1����M��y����E����   �e���M�a���ËT$�B�J�3���������������M����J����T$�B��J�3��������������hh�h�   hP��E�P�G�����ËT$�B��J�3������x������M��������T$�B��J�3��l����T��r����M��j����M��Ҫ���T$�BЋJ�3��A����0��G���������̍M��8����T$�BЋJ�3�������������M������T$�B�J�3�������d�������E����   �e���M�2���ÍM��)����T$�B�J�3������@������M������M�������T$�BԋJ�3������������M������M��ө���T$�B��J�3��b�������h����M��`����M�騩���T$�B��J�3��7����Ԫ�=����M��5����M��}����T$�B؋J�3�������������M��z����T$�B�J�3���������������M��W����T$�B�J�3�������h�������M��4����M��,����T$�B܋J�3������D������M���^���M���^���M�������T$�B��J�3��h���� ��n����M��֨���T$�B�J�3��E�������K����M��s^���T$�B��J�3��"����ة�(����M�� ����M��h����M��`����M��X����T$�B؋J�3���������������M�������T$�B�J�3���������������M�������T$�B�J�3������l������M������T$�B�J�3��~����H������M��|����M��ħ���T$�B؋J�3��S����$��Y����M��Q����M�陧���T$�B؋J�3��(���� ��.����M��V5���T$�B��J�3������ܨ�����M��s����T$�B��J�3���������������M��P����T$�B��J�3��������������M��-����T$�B�J�3������p������M��
����T$�B�J�3��y����L������M������E����   �e���M�Ϧ��ËT$�B�J�3��=����(��C����EЃ��   �e���M雦��ÍM�钦���M�銦���T$�BȋJ�3��������������M��g����M��_����M��W����M��O����M�������M��?����T$�B��J�3������������M������T$�B��J�3�������������M�������M������M������M��q����T$�B��J�3��P�������V����M��N����M��F����T$�B��J�3��%����t��+����M��#����T$�B�J�3������P������M��p����M��h����M��`����T$�BȋJ�3�������,�������M��=����T$�B��J�3������������̋E����   �e���M����ËT$�B��J�3��v����4��|��������������̍M�ؤ���T$�B��J�3��G����L��M���������������̍M��8����E܃��   �e���M� ���ËT$�B�J�3������� ��������̍M��(Z���Eԃ��   �e���M�Z��ËT$�B��J�3���������������̍M������M������E����   �e���M�ȣ��ËT$�BċJ�3��v�������|��������������̋M��أ���T$�B��J�3��G����\��M����M�鵣���T$�B��J�3��$����8��*����M�钣���T$�B��J�3������������M��o����T$�B��J�3��������������M��L����T$�B��J�3������̰������M��)����E����   �e���M����ËT$�B�J�3�������������M��X���M�����Eԃ��   �e���M�X��ÍM��Ģ���T$�B؋J�3��3�������9����M��aX���M院���Eԃ��   �e���M�AX��ÍM��x����T$�B؋J�3�������`�������M��X���Eԃ��   �e���M�=���ÍM��4����T$�B��J�3������<������M�����E����   �e���M�W��ËT$�B��J�3��g������m����M��ա���E����   �e���M齡��ËT$�B�J�3��+�������1����M�陡���T$�B�J�3������Я�����M��v����T$�B�J�3���������������M��S����T$�B�J�3���������������M���V���M�(����Eԃ��   �e���M��V��ÍM������T$�B؋J�3��v����d��|����M��V���M�ܠ���Eԃ��   �e���M�V��ÍM�黠���T$�B؋J�3��*����@��0����M�阠���E����   �e���M造��ËT$�B�J�3��������������M��V���M��T����T$�B��J�3���������������M���U���M�)����Eԃ��   �e���M��U��ÍM������T$�B؋J�3��w����Ԯ�}����M��U���M�ݟ���Eԃ��   �e���M�U��ÍM�鼟���T$�B؋J�3��+�������1����E����   �e���M��IU��ÍM�速���E����   �e���M��(U��ËM�_����E����   �e���M�U��ÍM��>����M��6����T$�B��J�3�������������M���T���M�����Eԃ��   �e���M�T��ÍM������T$�B؋J�3��Y����h��_����M��Ǟ���E����   �e���M鯞��ËT$�B�J�3������D��#�����̍M���{���E���   �e���M��{��ËT$�B��J�3�������d�������M��{���E���   �e���M�{��ËT$�B��J�3������@������M��{���E܃��   �e���M�h{��ËT$�B�J�3��f������l����E����   �e���M�ĝ��ÍM�黝���T$�B�J�3��*�������0����E���t�e���M錝��ËT$�B��J�3�������H�� ����M��h����M��`����T$�B��J�3�������$�������M��=����E����   �e���M�%���ËT$�B�J�3������ ������M������E����   �e���M����ËT$�B�J�3��W����ܵ�]����E���t�e���M�yR��ËT$�B��J�3��'�������-����E���t�e���M����ËT$�B��J�3���������������M��e����E����   �e���M�M���ËT$�B�J�3������p�������M��)����E����   �e���M����ËT$�B�J�3������L������M��Q���Eԃ�t�e���M�ٛ��ËT$�B��J�3��G����(��M����M�镛���E����   �e���M�}���ËT$�B�J�3������������M��	����M��Q����Ẽ��   �e���M����ËT$�BԋJ�3��������������M��5����E����   �e���M����ËT$�B�J�3�������������M��ٚ���E����   �e���M�����ËT$�B�J�3��O�������U����M��M����T$�B܋J�3��,����t��2����Ẽ��   �e���M銚��ÍM������M��Y����T$�BЋJ�3�������P�������Ẽ��   �e���M�F���ÍM��͹���M������T$�BЋJ�3������,������M�颹���M������T$�B؋J�3��y����������M��w����M�鿙���T$�B؋J�3��N������T����M��L����E܃�t�e���M�8���ËT$�B�J�3�����������������������̍M�8O���T$�B��J�3�������t������������������̍M��ظ���E܃�t�e���M�ĸ��ËT$�B�J�3������м�����M�頸���E܃�t�e���M錸��ËT$�B�J�3��j�������p����M�鸘���M��@v���T$�BԋJ�3��?�������E����M�鍘���M��v���T$�B؋J�3������d������M��b����M���u���Ẽ��   �e���M�"N��ËT$�BЋJ�3�������@�������M������M��u���Ẽ��   �e���M��M��ËT$�BЋJ�3������������M��ڗ���M��bu���T$�B؋J�3��a�������g����M�鯗���M��7u���T$�B؋J�3��6����Ի�<����M�鄗���M��u���T$�B̋J�3�������������M��Y����M��t���T$�B��J�3���������������M��.����M��t���T$�BԋJ�3������h������M������M��t���T$�B؋J�3������D������M��ؖ���M��`t���T$�BԋJ�3��_���� ��e����M�魖���M��5t���T$�B؋J�3��4�������:����M�邖���M��
t���T$�BԋJ�3��	����غ�����M��W����M���s���T$�B؋J�3���������������M��,����M��s���T$�BԋJ�3�������������M������M��s���T$�B؋J�3������l������M��֕���M��^s���T$�BԋJ�3��]����H��c����M�髕���M��3s���T$�B؋J�3��2����$��8����M�逕���M��s���T$�BԋJ�3������ ������M��U����M���r���T$�B؋J�3�������ܹ������M��*����M��r���T$�BԋJ�3�������������M�������M��r���T$�B؋J�3�������������M��Ԕ���M��\r���T$�BԋJ�3��[����p��a����M�驔���M��1r���T$�B؋J�3��0����L��6����M��~����M��r���T$�BԋJ�3������(������M��S����M���q���T$�B؋J�3��������������M��س���M�������T$�BċJ�3������������M��͂���M������T$�B܋J�3�������������M�颂���M��j����T$�B܋J�3��Y�������_������������������hЃ����Y����̃=� uK����t� �Q�@<�@�Ѓ���    V�5���t���0I��V�
�������    ^�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           �� l� R� 6� "� � � ��     ھ � �� � � "� *� 4� ¾ P� Z� h� ~� �� �� Ŀ � �� �� �� �� �� p� B� d�         ��        f\�_            �������N���������������C-DT�!	@-DT�!�?tristate-undef.tif  tristate-on.tif tristate-off.tif    tristate-multiple.png   src/TriStateGui.cpp src/TriStateGui.cpp Tristate    �������N    ���������������C-DT�!	@-DT�!�?|�@ �S �S � �S �S �   PT `T pT ��� � P �d  �d �d �d Ц � @ p `� p� ��   � �� Ч � � P�� � ` � � �< � src/TriStateGui.cpp TRISTATE    ../../resource/_api/c4d_resource.cpp    ../../resource/_api/c4d_resource.cpp    #   #   #   #   #   #   #   #   #   #   M_EDITOR    M_EDITOR    ���6 res �������N    ���������������C-DT�!	@-DT�!�?�������N���������������C-DT�!	@-DT�!�?../../resource/_api/c4d_basebitmap.cpp  ../../resource/_api/c4d_basebitmap.cpp  ../../resource/_api/c4d_basebitmap.cpp  ../../resource/_api/c4d_basebitmap.cpp  ../../resource/_api/c4d_basebitmap.cpp  �������N���������������C-DT�!	@-DT�!�?p:\applications\maxon\cinema 4d r14.041\resource\_api\c4d_misc/datastructures/basearray.h       ~   Progress Thread 0%  ../../resource/_api/c4d_gui.cpp ../../resource/_api/c4d_gui.cpp %   ../../resource/_api/c4d_gui.cpp ../../resource/_api/c4d_gui.cpp ../../resource/_api/c4d_gui.cpp ../../resource/_api/c4d_gui.cpp ../../resource/_api/c4d_gui.cpp �������N    ���������������C-DT�!	@-DT�!�?ܛ�� �S �S �S �S �S  T @T PT `T pT țp� `d pd �d �d �d �d �d �d �p� `d pd �d �d �d �d �d �� ��p� `d pd �d �d �d �d �d p� <�p� `d pd �d �d �d �d �d Ц 0� @� P� `� p� �� �� �� �� Ч � �       �?-DT�!	@      Y@     �f@     @�@�������������../../resource/_api/c4d_file.cpp    ../../resource/_api/c4d_file.cpp    �������N���������������C-DT�!	@-DT�!�?%s     p:\applications\maxon\cinema 4d r14.041\resource\_api\c4d_general.h ../../resource/_api/c4d_basetime.cpp    ../../resource/_api/c4d_basetime.cpp    ../../resource/_api/c4d_basetime.cpp        ����MbP?      �?   ����A  4&�kC �Ngm��C  4&�k�        ��������������       �       �P��*+�[�[    �������N���������������C-DT�!	@-DT�!�?../../resource/_api/c4d_pmain.cpp   ../../resource/_api/c4d_pmain.cpp   ��\    X���    H                                                           P����              x�����    �       ����    @   h�0�        ����    @   ��           ̙��    H�       ����    @   �            �ԙ�H�    d�       ����    @   ,�           <��H�    |�        ����    @   d�           t�H�                ����           ����Ț    ��       ����    @   ����        ����    @   �           ��Ț                ���            �4�ԙ�H�    ��       ����    @   �            ��d�           t�������    ��       ����    @   d�            0���            d�,�            |�d�            ���            ��           � �H�    �       ����    @   �            H��             �d�           t�|�     �        ����    @   d�            8���           ��Ĝ    8�        ����    @   ���e @f kf �f g Cg hg �g �g (h Xh �h �h i pi �i !j vj �j �j Vk �k �k  l &l ]l �l �l �l �l 7m bm �m �m �m n )n Tn �n �n �n o +o No qo �o �o �o p 0p Sp vp �p �p Aq dq �q �q �q  r Cr yr �r �r 1s ys �s �s �s t 4t pt �t u Lu �u �u �u 
v -v yv �v w ,w xw �w Jx �x �x y My �y �y �y  z \z �z �z �z 4{ p{ �{ �{ (| d| �| �| } K} v} �} �} ~ M~ �~ �~ �~  c � � � � :� e� �� �� � � <� g� �� �� � � >� i� �� �� � � @� k� ��                 ����0g    ;g"�   0�                       �����f����[f    cf����0f    8f"�
   �                       "�   d�                       "�   l�                       "�   |�                       �����f    �f�����f   �f�����f   �f�����f   �f�����f����g���� h"�   l�                       �����g    �g   �g"�   ��                       ����`g"�   Ԡ                       �����g    �g"�    �                       ����sh����Ph����<j����Dj   ]j�����i�����i   j�����h    �h   �h�����h    �h   �h   i"�   D�                       "�   \�                       "�   ��                       "�   ̢                       "�   ��                       "�   t�                       "�   4�                       "�   <�                       ����Gi    7i   ?i   `i   hi�����i    �i   �i   �i   �i   �i�����j    �j"�   $�                       �����j    �j"�   X�                       "�   ��                       ���� k    +k   6k   >k   Fk   Nk����xl����Al����l�����k�����l�����l�����k    �k�����k    �k"�    �                       "�   �                       "�   �                       "�   �                       "�   �                       "�   ��                       "�    �                       ����`r"�   ,�                       ����;r�����q����\q����np����Kp����(p����p�����o����io����Fo����#o�����n�����n����!n�����m�����l�����l�����q�����q�����p    �p�����o    �o�����o    �o����Dn    Ln�����m    �m�����m    �m����}m    �m����Rm    Zm����m    /m����r    r   r�����p    �p    �p����on    wn   n����q    �q   �q�����q�����n    �n    �n     o"�   X�                       "�   ��                       "�   `�                       "�   �                       "�   Ȧ                       "�   h�                       "�   ��                       "�   ��                       "�   �                       "�   p�                       "�   x�                       "�   ��                       "�   ��                       "�   ��                       "�    �                       "�   �                       "�   ��                       "�   ��                       "�   ��                       "�   �                       "�   ��                       "�   ��                       "�   ��                       "�    �                       "�   ��                       "�   ȥ                       "�   0�                       "�   @�                       "�   P�                       "�   `�                       "�   p�                       "�   Х                       "�   إ                       ����q����q����!q����)q����1q   9q����s    s"�   ܫ                       �����r    �r"�   �                       �����r"�   D�                       ����`s    Xs    Ps"�   p�                       ����%v����v�����u����,t����	t�����s�����s�����s�����x    �x����w����$w�����v    �v�����u    �u����ou    gu����Wt    Ot����+u    #u    Du����ux    ex   mx    �x�����w    �w   �w    �w����Ww    Gw   Ow    pw�����v    �v   �v    �v����Xv    Hv   Pv    qv�����t    �t   �t     u�����t    �t   �t    �t"�   �                       "�   d�                       "�   ��                       "�   ��                       "�   ��                       "�   ��                       "�   �                       "�   ĭ                       "�   �                       "�   ��                       "�   ��                       "�   ��                       "�   �                       "�   ,�                       "�   L�                       "�   �                       "�   $�                       "�   <�                       "�   Ĭ                       "�   ̬                       "�   Ԭ                       "�   ܬ                       "�   �                       ����!x    �w   �w    x   x   :x    Bx�����y    �y����py    hy����4y    ,y�����x    �x"�   ��                       "�   ȱ                       "�   ر                       "�   �                       �����|�����z�����z�����y�����}    �}�����}    �}����f}    n}�����|    |����K|    C|�����{    �{�����{    �{����W{    O{����{    {����z    wz����Cz    ;z����"}    ;}   C}�����|    �|   �|����z    z����z����|    �{   |    |"�   ��                       "�   ��                       "�   Ȳ                       "�   X�                       "�   p�                       "�   ��                       "�   ز                       "�   �                       "�   ��                       "�   ��                       "�   �                       "�   �                       "�   (�                       "�   ��                       "�   ��                       "�   8�                       "�   H�                       "�   ��                       "�   ��                       ���� ~"�   l�                       ������    ������[�    c�����0�    8������    �����ڂ    �������    ��������    ������Y�    a�����.�    6������    �����؁    ��������    ��������    ������W�    _�����,�    4������    	�����ր    ހ������    ��������    ������U�    ]�����*�    2������    ������    ������    �����~    ������~    �~�����~    �~����p~    h~����8~    0~����J    :   B����    �~   �~"�   ��                       "�   ��                       "�   ��                       "�   ȶ                       "�   ض                       "�   �                       "�   ��                       "�   �                       "�   �                       "�   (�                       "�   8�                       "�   H�                       "�   X�                       "�   h�                       "�   x�                       "�   ��                       "�   ��                       "�   ��                       "�   ��                       "�   ȷ                       "�   ط                       "�   �                       "�   ��                       "�   �                       "�   �                       "�   h�                       "�   ��                       "�   (�                       "�   8�                       "�   H�                       "�   X�                           ����    ����    ����    �_    �_�_����    ����    ����    �`    ����    ����    ����    �b    ����    ����    �����b�b    ����    ����    ����	dd��         �� $� ؽ         ��  �                     �� l� R� 6� "� � � ��     ھ � �� � � "� *� 4� ¾ P� Z� h� ~� �� �� Ŀ � �� �� �� �� �� p� B� d�     1_purecall x__CxxFrameHandler3  ,memset  �free  malloc  �floor Q_CIfmod MSVCR110.dll  p ??1type_info@@UAE@XZ  s__CppXcptFilter _amsg_exit  �_malloc_crt �_initterm �_initterm_e |_lock �_unlock +_calloc_crt �__dllonexit "_onexit 
_vsnprintf  K_crt_debugger_hook  �__crtUnhandledException �__crtTerminateProcess ;?terminate@@YAXXZ �__clean_type_info_names_internal  p_except_handler4_common <EncodePointer DecodePointer �IsDebuggerPresent �IsProcessorFeaturePresent <QueryPerformanceCounter $GetCurrentProcessId (GetCurrentThreadId  �GetSystemTimeAsFileTime KERNEL32.dll      ��R    ��          �� �� �� 0T �   tristategui.cdl c4d_main                                                                                                                                                                                                                                                      
   
            �    .?AVCustomGuiData@@ �    .?AVBaseData@@  �    .?AViCustomGui@@    �    .?AVSubDialog@@ �    .?AVGeDialog@@  �    .?AVTriStateUA@@    �    .?AVGeUserArea@@    �    .?AVTriStateGui@@   �    .?AVTriStateData@@  �    .?AVGeModalDialog@@ �    .?AVC4DThread@@ �    .?AVtype_info@@ N�@���D        ����                                                                                                                                                               �   -0S0c0�0�0�0�0C1S1�1�1�12
2c2q2�2�2�233A3S3f3�3�3�3�3 4U4[4u4�4�4�4�45!545�5�5�5�5�5�56-6a6k6u66�6�6�67A7a7�7�7�7c8r8�8�8�8�9::::$:3:T:Z:`:f:x:|:�:�:�:�:�:3;Q;�;�;�;�;�;�;<<*<H<t<�<�<
=/=�=�=�=�=8>Q>�>�>?*?@?E?i?�?�?�?       0060e0�0�0�0S1a1}1�1+2S2�2�23333D3_3i3u3�3�3�3�3�3�34(4B4�4�4�4�455/595E5X5o5�5�5�5�5�5�56W6t6�6�6�6�6�67,7>7R7�7�7�7�7�7�7�78,8?8J8n8�8�8�899)949X9r9�9�9�9�9�9:*:L:i:{:�:�:�:�:	;;(;?;R;l;;�;�;�;�;'<D<V<i<t<�<�<�<�<=!=,=P=j=�=�=�=�=�=�=>9>V>h>|>�>�>D?Y?|?�?�?�?   0  �    00010�0�01>1g1�1�1�122"292�2�23@3i3�3�3444$464A4[4s4�4�4�4�4�4"525Q5a5s5�5�5�566!616A6Q6a6q6�6�6�6�6�67!7Q7q7�7�7�7�78818N8q8�9�9�9�9�9�9�9�9�9�9�9�9�9::::�:�:�:
;;�;(=0=8=@=H=P=�=�=�=>1>`>�>�>�>�>?$?B?[?u?�?�?�?   @  �   0!0A0Q0a0q0�0�0�0�0!1E1q1�1�1�1�1�1�112E2e2�2�2�23A3T3i3�3�3�34!4A4a4�4�4�4�4�45A5\5�5�5�56/6D6N6�677o7�7�7�78!818�8�8�9�9�9:c:q:�:7;<;�;�<=!=1=Q=a=#?5?�?�?�?�?   P  �   �0�0C2�2�223Y3`3�3�3r4�4 595U5o5+6c6s6�6�67Q7q7�7�7�7�7858e8�8�8�8�89 949X9l9�9�9�9�9:1:Q:r:�:�:�:�:�:;*;K;_;s;�;�;�;�;�;%<Q<w<�<�<=E==�=>1>U>�>�>�>�>!?A?e?�?�?�?   `  �   0E0c0t0�0�01*1U1�1�1�1242k2�2�2�2[3�3�3�344484A4�45M56<6{6�6�6�67?7Z7�7�7�78A8h8�8�8�8(9h9�9�9�9:3:M:g:�:�:�:�:;i;y;�;�;�;<(<K<�<�<�<�<=�=�=�=�=h>�>�>?�?�?   p  �   %0�0�0�0�0�0�0.1G1�1�1�1�12B2X2�2�23@3�3�3(4n4�4�45:5W5�5�56,6D6�6�6�6�687a7�7�7�8*9Z9b9j9�9�9%:�:�:;#;7;�;�;�;�;B<�<�<�<g=�=�=>->e>�>�>�>A?m?�?�?�?   �  �   00E0a0�0�0�0Z1�1�133;3K3g3�3�4�4�45I5i5�5�56a6�6�6�6-7U7�7�788?8�8�8?9�9�9/::�:;o;�;<_<�<�<O=�=�=/>>�>?h?�?   �  �   	0*0�0�01M1�1�12A2q2�2�23=3q3�3�3�3K4�4�4�4
555e5~5�5�56Y6�6�6�6+7k7�7�7�7!8Q8�8�8�89A9�9�9�9�9:&:�:�:�:;/;I;�;<;<s<�<�<�<==-=A=q=�=�=�=�=>c>s>�>�>�>�>V?[?`?z?�?�?�?�?   �  �   d0�0�0%1�12|2�2�2�2�2�2�2�2�2�2�34444 4$4(4,404555*5H5Q5q5�566*6/686^6f6�6�6�6S8b8�8�8�89�9�9�9#:3:l:�:�:;;#;4;R;n;�;�;�;�; <<M<u<�<�<�<�<�<==3=J=l=�=�=�=>#>5>g>�>�>�>�>?3?s?�?�?�?   �  �   0:00�0�0�031D11�1�1�1�132D2X2j2}2�2�233I3f3�3�3�3 44S4d4x4�4%5W5�5�536�6�6�6�6�6�67;7Y7u7�7�7�7�7>8T8�8�89<9�9�9�9�9�9:%:<:L:i:�:�:�:�:;`;s;�;�;B<a<�<V=u=�=�=�>�>�?�? �  �   f0�0�0�1�1�122:2x2�2�2�2C4P4y4�4�4�45 5s5�5�56626G6a6q6�8�899h9�9W:^:e:l:s:z:�:�:�:�:�:�:�:;!;5;S;a;y;�;�;�;�;�;<C<Q<i<w<�<�<�<�<�<=C=Q=i==�=�=�=>>.>D>^>n>�>�>�>�>?.?A?X?s?�?�?�?�?   �    0!080S0�0�0�0�011A1Q1q1�1�1�1�12!212S2a2{2�2�2�23!3A3c3t3�3�3�3�34!414A4Q4a4�4�4�4�4�4�4�455!515A5Q5a5q5�5�5�5�5�526s6�6�6�6�6�6 757�7�7�78A8[8r8�8�8�8�8	9 9q9�9�9�9�9�9A:Q:a:q:�:�:�:�:�:;#;3;f;�;�;�;�;�;.<B<�<�<�<=&=F=�=�=�=�=>0>N>l>�>�>�>?B?b?�?�?�?   �  p  00!010Q0q0�0�0�0�0�0�0�0�01#1=1P1g1�1�1�122#242N2c2}2�2�2�23323G3a3q3�3�3�3�344!414A4Q4a4q4�4�4�4�45!515A5Q5a5q5�5�5�5�5�5�5�566A6Q6a6q6�6�6�6�6�6�6�6�677!717A7Q7a7q7�7�7�7�7�7�7�7!8A8Q8a8q8�8�8�8�8�8�8�8�899A9Q9a9q9�9�9�9�9�9�9�9�9:%:F:r:�:�:�:;;!;1;A;Q;c;t;�;�;�;�;�;<3<D<^<v<�<�<�<�<3=E=`=�=�=�=�=�=>+>Y>t>�>�>�>�>?'?>?Y?�?�?�?�?�?�?   �  �   0(080q0�0�0�0�0�01A1q1R2�2�2�23b3�3�3�34B4j4�4�4�4"5R5�5�5�5�526r6�6�6�6!7l7�7�7�78a8�8�8�8�899:9`9�9�9�9#:3:E:�:�:;a;�;�;"<b<�<�<=B=�=�=�=B>r>�>�>2?r?�?�?     0B0�0�0131C1W1�1�162�2�23R3�3�3"4b4�4�4#545F5i5�5�5�5616Q6q6�6�6�67757Q7q7�7�7�78%8A8e8�8�8�8�899#919K9f9�9�9�9�9�9�9::%:Q:c:r:�:�:�:�:�:�:1;A;S;d;~;�;�;�;<<.<F<`<p<�<�<�<�<�<==!=1=A=Q=a=q=�=�=�=�=�=�=�=�=>a>q>�>�>�>�>�>�>1?A?Q?�?�?�?      00!010A0Q0a0q0�0�0�0�0�0�0�0
1$141s1�1�1�1�1�1!212D2t2�2�2�2�233!313A3S3b3�3�3�344'4O4d4i4�4�4�4$5U5�5�5�56%6Q6a6�6�6�6�67S7c7�7�7 8A8Q8a8s8�8�8�8�8�839C9e9�9�9�9::::\:�:�:�:�:;I;�;�;�;�;<$<><R<�<�<�<�<�<S=c=u=�=�=�=C>S>e>�>�>�>1?A?Q?l?�?�?�?�?�?�?�?        00!010A0Q0a0s0�0�011!111A1Q1a1q1�1�1�1�1�1�1�1�122C2Q2c2�2!3Q3w3�3�3�3+474�4�45+5<5G5a5�5�5�5�56(6-6B6]6�6�6�6�6�6�6�6
7�7�7�7�7�7�7�78H8h8�8�8�89999C9Y9�9�9:!:A:a:�:�:�:�:�:�:!;A;a;w;�;�;�;<<1<A<c<r<�<�<=1=Q=q=�=�=�=�=!>A>a>�>�>�>�>�>�>??!?1?A?Q?q?�?�?�?�?�?   0 �   010S0b0�0�0�0y1�1�1�1[2�2�283[3�3�3H4k4�4�4�4W5�5�5�576s6�67,7s7�7�738D8�8�8#939�9�9�9v:�:�:�:;#;7;�;�;<�<�<�<�<#=3=G=�=>A>�>�>?1?O?m?�?�?�?   @ �   W0�0�0&1A1_1}1�1�1�1g2�2�293T3�3�34S4d4�455=5�5�5�5'6c6t6�67S7c7�78$8�8�899�9�9:%:Q:q:�:�:�:�:�:f;�;�;�;�;<'<F<c<q<�<�<=1=Q=q=�=�=�=�=>5>e>�>�>�>�>�>??!?1?A?Q?p?u?z??�?�?�?�?�?   P <  00A0W0}0�0�0�0�0#131}1�1�1C2S2�2�2
3a3q3�3�34B4N4T4�4�4�4�455 5$5(5,505K5T5�5�5�5�566!616A6a6�6�6�6�6707q7�7�7�7�718Q8q8�8�8�8�8�8�8�899!919A9Q9a9q9�9�9�9�9�9�9�9�9!:1:Q:q:�:�:�:�:;4;J;\;�;�;�;�;�;<<<*<n<x<}<�<�<�<�<�<�<==#=6=<=V=b=k=u={=�=�=�=�=�=�=�=>">5>:>@>T>Y>e>t>|>�>�>�>�>�>	?s?�?�?   `     000!0&0=0H0N0a0v0�0�0�0�01111+1c1i1o1u1{1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�122.272E2�2333�3�3�3�3�3�3x4�4�4�4�4�4�4555.535N5T5Y5q5�5�5�5�5�5�5 666666$6R6}6�6�6�67U7z7�7�7�78:8j8t8{8�8�8.9�9�93:�:�:;n;�;�;<8<B<L<o<�<�<�<=I=t=�=�=�=>;>f>�>�>�>?=?`?�?�?�?�? p �   0B0e0�0�01S1v1�1�1�122U2�2�23C3�3�3�3 4#4F4�4�45^5�5�5�56?6�6�67>7�7�7\8�8�8#9_9�9�9:2:n:�:�:
;F;�;�;�;:<v<�<�<=]=�=�=�=>_>�>�>�>1?u?�?�?�? � D   !0L0w0�0�0�0#1N1y1�1�1�1%2P2{2�2�2�2'3R3}3�3�3�3�3�3�344   � �  �0�0�0�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1 22222222 2$2(2,2�2�2�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5 66666666 6$6(6,6064686<6@6D6H6L6P6T6X6\6`6d6h6l6p6t6x6|6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�8�8�8�8�89999\9`9t9x9|9�9�9�9�9�9�9�9�9�9 ::::(:8:<:@:H:`:p:t:�:�:�:�:�:�:�:�:�:�:�:;;; ;$;(;,;4;L;\;`;p;t;x;|;�;�;�;�;�;�;�;�;�;�;�; <<<< <8<H<L<\<`<p<t<|<�<�<�<�<�<�<�<4?<?H?h?p?x?�?�?�?�?�? �    0 0(00080@0H0P0X0`0h0p0|0�0�0�0�0�0�011181@1H1P1X1`1h1p1x1�1�1�1�1�1�1�1�1�1 2D2h2�2�2�2�2�2�2�2�2 3333 3(303<3\3d3p3�3�3�3�3�3�3�3�3�3�3�34444$4,484\4�4�4�4�4505<5\5d5l5t5|5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�56666$6,646<6D6L6T6\6d6l6t6|6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�67747X7|7�7�7�7808T8x8�8�8�89,9P9t9�9�9�9:(:L:p:�:�:�: ;$;H;l;�;�;�;�;�;�;�;�;�;�;<<(<H<T<t<|<�<�<�<�<�<�<�<�<�<�<�<�< ==== =(=0=8=@=H=P=X=`=h=p=x=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�= >>>> >(>0>8>@>L>p>�>�>�> ?$?H?l?�?�?�?�?   � �   0D0h0�0�0�0�01@1d1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1 2$2H2l2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�23333$3,343<3D3L3T3\3d3l3t3|3�3�3�3�3�3�3�3�3�3�3444X4|4�4�4�4505T5x5�5�5�56,6P6p6|6�6�6�6�6�6�6�6�6�6�6�6�6�67777$7,747<7D7L7T7\7d7l7t7|7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�78888$8,848<8D8L8T8\8d8l8t8|8�8�8�8�8�8�8909T9x9�9�9�9:,:P:t:�:�:�:;(;L;p;�;�;�; <$<H<l<�<�<�<===8=X=t=x=�=�=   �     000H0d0|0�0�0�0�01 181                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                